// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    io_in,
    io_oeb,
    io_out,
    la_data_out);
 input wb_clk_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [63:0] la_data_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.alu_op[0] ;
 wire \as2650.alu_op[1] ;
 wire \as2650.alu_op[2] ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[10] ;
 wire \as2650.cycle[11] ;
 wire \as2650.cycle[12] ;
 wire \as2650.cycle[13] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.cycle[8] ;
 wire \as2650.cycle[9] ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ivec[0] ;
 wire \as2650.ivec[1] ;
 wire \as2650.ivec[2] ;
 wire \as2650.ivec[3] ;
 wire \as2650.ivec[4] ;
 wire \as2650.ivec[5] ;
 wire \as2650.ivec[6] ;
 wire \as2650.ivec[7] ;
 wire \as2650.last_intr ;
 wire \as2650.prefixed ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[10][0] ;
 wire \as2650.stack[10][10] ;
 wire \as2650.stack[10][11] ;
 wire \as2650.stack[10][12] ;
 wire \as2650.stack[10][13] ;
 wire \as2650.stack[10][14] ;
 wire \as2650.stack[10][1] ;
 wire \as2650.stack[10][2] ;
 wire \as2650.stack[10][3] ;
 wire \as2650.stack[10][4] ;
 wire \as2650.stack[10][5] ;
 wire \as2650.stack[10][6] ;
 wire \as2650.stack[10][7] ;
 wire \as2650.stack[10][8] ;
 wire \as2650.stack[10][9] ;
 wire \as2650.stack[11][0] ;
 wire \as2650.stack[11][10] ;
 wire \as2650.stack[11][11] ;
 wire \as2650.stack[11][12] ;
 wire \as2650.stack[11][13] ;
 wire \as2650.stack[11][14] ;
 wire \as2650.stack[11][1] ;
 wire \as2650.stack[11][2] ;
 wire \as2650.stack[11][3] ;
 wire \as2650.stack[11][4] ;
 wire \as2650.stack[11][5] ;
 wire \as2650.stack[11][6] ;
 wire \as2650.stack[11][7] ;
 wire \as2650.stack[11][8] ;
 wire \as2650.stack[11][9] ;
 wire \as2650.stack[12][0] ;
 wire \as2650.stack[12][10] ;
 wire \as2650.stack[12][11] ;
 wire \as2650.stack[12][12] ;
 wire \as2650.stack[12][13] ;
 wire \as2650.stack[12][14] ;
 wire \as2650.stack[12][1] ;
 wire \as2650.stack[12][2] ;
 wire \as2650.stack[12][3] ;
 wire \as2650.stack[12][4] ;
 wire \as2650.stack[12][5] ;
 wire \as2650.stack[12][6] ;
 wire \as2650.stack[12][7] ;
 wire \as2650.stack[12][8] ;
 wire \as2650.stack[12][9] ;
 wire \as2650.stack[13][0] ;
 wire \as2650.stack[13][10] ;
 wire \as2650.stack[13][11] ;
 wire \as2650.stack[13][12] ;
 wire \as2650.stack[13][13] ;
 wire \as2650.stack[13][14] ;
 wire \as2650.stack[13][1] ;
 wire \as2650.stack[13][2] ;
 wire \as2650.stack[13][3] ;
 wire \as2650.stack[13][4] ;
 wire \as2650.stack[13][5] ;
 wire \as2650.stack[13][6] ;
 wire \as2650.stack[13][7] ;
 wire \as2650.stack[13][8] ;
 wire \as2650.stack[13][9] ;
 wire \as2650.stack[14][0] ;
 wire \as2650.stack[14][10] ;
 wire \as2650.stack[14][11] ;
 wire \as2650.stack[14][12] ;
 wire \as2650.stack[14][13] ;
 wire \as2650.stack[14][14] ;
 wire \as2650.stack[14][1] ;
 wire \as2650.stack[14][2] ;
 wire \as2650.stack[14][3] ;
 wire \as2650.stack[14][4] ;
 wire \as2650.stack[14][5] ;
 wire \as2650.stack[14][6] ;
 wire \as2650.stack[14][7] ;
 wire \as2650.stack[14][8] ;
 wire \as2650.stack[14][9] ;
 wire \as2650.stack[15][0] ;
 wire \as2650.stack[15][10] ;
 wire \as2650.stack[15][11] ;
 wire \as2650.stack[15][12] ;
 wire \as2650.stack[15][13] ;
 wire \as2650.stack[15][14] ;
 wire \as2650.stack[15][1] ;
 wire \as2650.stack[15][2] ;
 wire \as2650.stack[15][3] ;
 wire \as2650.stack[15][4] ;
 wire \as2650.stack[15][5] ;
 wire \as2650.stack[15][6] ;
 wire \as2650.stack[15][7] ;
 wire \as2650.stack[15][8] ;
 wire \as2650.stack[15][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \as2650.stack[8][0] ;
 wire \as2650.stack[8][10] ;
 wire \as2650.stack[8][11] ;
 wire \as2650.stack[8][12] ;
 wire \as2650.stack[8][13] ;
 wire \as2650.stack[8][14] ;
 wire \as2650.stack[8][1] ;
 wire \as2650.stack[8][2] ;
 wire \as2650.stack[8][3] ;
 wire \as2650.stack[8][4] ;
 wire \as2650.stack[8][5] ;
 wire \as2650.stack[8][6] ;
 wire \as2650.stack[8][7] ;
 wire \as2650.stack[8][8] ;
 wire \as2650.stack[8][9] ;
 wire \as2650.stack[9][0] ;
 wire \as2650.stack[9][10] ;
 wire \as2650.stack[9][11] ;
 wire \as2650.stack[9][12] ;
 wire \as2650.stack[9][13] ;
 wire \as2650.stack[9][14] ;
 wire \as2650.stack[9][1] ;
 wire \as2650.stack[9][2] ;
 wire \as2650.stack[9][3] ;
 wire \as2650.stack[9][4] ;
 wire \as2650.stack[9][5] ;
 wire \as2650.stack[9][6] ;
 wire \as2650.stack[9][7] ;
 wire \as2650.stack[9][8] ;
 wire \as2650.stack[9][9] ;
 wire net142;
 wire net147;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net143;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net144;
 wire net112;
 wire net113;
 wire net114;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net145;
 wire net146;
 wire net115;
 wire net120;
 wire net116;
 wire net117;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net118;
 wire net119;
 wire net153;
 wire net126;
 wire net154;
 wire net127;
 wire net155;
 wire net128;
 wire net156;
 wire net129;
 wire net157;
 wire net130;
 wire net158;
 wire net131;
 wire net159;
 wire net132;
 wire net160;
 wire net133;
 wire net134;
 wire net161;
 wire net135;
 wire net162;
 wire net136;
 wire net163;
 wire net137;
 wire net164;
 wire net138;
 wire net165;
 wire net139;
 wire net166;
 wire net140;
 wire net167;
 wire net141;
 wire clknet_leaf_0_wb_clk_i;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_leaf_130_wb_clk_i;
 wire clknet_leaf_131_wb_clk_i;
 wire clknet_leaf_132_wb_clk_i;
 wire clknet_leaf_133_wb_clk_i;
 wire clknet_leaf_134_wb_clk_i;
 wire clknet_leaf_135_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire clknet_opt_2_0_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05815_ (.I(\as2650.cycle[6] ),
    .ZN(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05816_ (.I(_05669_),
    .Z(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05817_ (.I(_05670_),
    .Z(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05818_ (.I(_05671_),
    .Z(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05819_ (.I(_05672_),
    .Z(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05820_ (.I(_05673_),
    .Z(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05821_ (.I(net5),
    .Z(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05822_ (.I(_05675_),
    .Z(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05823_ (.I(_05676_),
    .Z(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05824_ (.I(_05677_),
    .Z(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05825_ (.I(\as2650.ins_reg[4] ),
    .ZN(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05826_ (.I(_05679_),
    .Z(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05827_ (.I(_05680_),
    .Z(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05828_ (.I(net94),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05829_ (.I(\as2650.ins_reg[0] ),
    .Z(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05830_ (.I(_05683_),
    .Z(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05831_ (.I(_05684_),
    .Z(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05832_ (.A1(_05682_),
    .A2(_05685_),
    .Z(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05833_ (.I(net54),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05834_ (.I(\as2650.ins_reg[1] ),
    .Z(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05835_ (.A1(_05687_),
    .A2(_05688_),
    .Z(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05836_ (.A1(_05686_),
    .A2(_05689_),
    .ZN(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05837_ (.I(\as2650.alu_op[2] ),
    .Z(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05838_ (.I(\as2650.alu_op[1] ),
    .Z(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05839_ (.I(_05692_),
    .Z(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05840_ (.I(_05693_),
    .ZN(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05841_ (.A1(_05691_),
    .A2(_05694_),
    .ZN(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05842_ (.I(_05688_),
    .Z(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05843_ (.A1(_05696_),
    .A2(_05685_),
    .ZN(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05844_ (.A1(_05697_),
    .A2(_05690_),
    .ZN(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05845_ (.I(\as2650.ins_reg[4] ),
    .Z(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05846_ (.I(_05699_),
    .Z(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05847_ (.A1(_05691_),
    .A2(_05693_),
    .ZN(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05848_ (.A1(_05700_),
    .A2(_05701_),
    .ZN(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _05849_ (.A1(_05681_),
    .A2(_05690_),
    .A3(_05695_),
    .B1(_05698_),
    .B2(_05702_),
    .ZN(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05850_ (.I(_05700_),
    .Z(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05851_ (.I(\as2650.ins_reg[0] ),
    .Z(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05852_ (.A1(\as2650.ins_reg[1] ),
    .A2(_05705_),
    .Z(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05853_ (.I(_05706_),
    .Z(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05854_ (.I(_05707_),
    .Z(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05855_ (.I(net51),
    .Z(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05856_ (.I(_05709_),
    .Z(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05857_ (.I(_05710_),
    .Z(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05858_ (.I(_05711_),
    .Z(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05859_ (.I(_05712_),
    .Z(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05860_ (.I(_05713_),
    .Z(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05861_ (.I0(\as2650.r123[1][7] ),
    .I1(\as2650.r123[0][7] ),
    .I2(\as2650.r123_2[1][7] ),
    .I3(\as2650.r123_2[0][7] ),
    .S0(_05685_),
    .S1(_05714_),
    .Z(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05862_ (.A1(_05708_),
    .A2(_05715_),
    .ZN(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05863_ (.A1(\as2650.ins_reg[1] ),
    .A2(_05705_),
    .Z(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05864_ (.I(_05717_),
    .Z(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05865_ (.I(_05718_),
    .Z(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05866_ (.I(_05719_),
    .Z(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05867_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_05713_),
    .Z(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05868_ (.A1(_05720_),
    .A2(_05721_),
    .ZN(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05869_ (.I(\as2650.r0[7] ),
    .Z(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05870_ (.I(_05723_),
    .Z(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05871_ (.A1(_05688_),
    .A2(_05683_),
    .ZN(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05872_ (.I(_05725_),
    .Z(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05873_ (.I(_05726_),
    .Z(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05874_ (.I(_05727_),
    .Z(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05875_ (.A1(_05724_),
    .A2(_05728_),
    .ZN(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05876_ (.A1(_05716_),
    .A2(_05722_),
    .A3(_05729_),
    .ZN(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05877_ (.I(\as2650.r0[5] ),
    .Z(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05878_ (.I(_05731_),
    .Z(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05879_ (.I(_05732_),
    .Z(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05880_ (.I(_05726_),
    .Z(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05881_ (.A1(_05733_),
    .A2(_05734_),
    .ZN(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05882_ (.I(_05712_),
    .Z(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05883_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_05736_),
    .Z(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05884_ (.I0(\as2650.r123[1][5] ),
    .I1(\as2650.r123[0][5] ),
    .I2(\as2650.r123_2[1][5] ),
    .I3(\as2650.r123_2[0][5] ),
    .S0(_05684_),
    .S1(_05736_),
    .Z(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05885_ (.I(_05707_),
    .Z(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05886_ (.A1(_05719_),
    .A2(_05737_),
    .B1(_05738_),
    .B2(_05739_),
    .ZN(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05887_ (.A1(_05735_),
    .A2(_05740_),
    .Z(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05888_ (.I(\as2650.r0[6] ),
    .Z(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05889_ (.I(_05742_),
    .Z(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05890_ (.A1(_05743_),
    .A2(_05727_),
    .ZN(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05891_ (.I(_05718_),
    .Z(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05892_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_05713_),
    .Z(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05893_ (.I0(\as2650.r123[1][6] ),
    .I1(\as2650.r123[0][6] ),
    .I2(\as2650.r123_2[1][6] ),
    .I3(\as2650.r123_2[0][6] ),
    .S0(_05684_),
    .S1(_05713_),
    .Z(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05894_ (.A1(_05745_),
    .A2(_05746_),
    .B1(_05747_),
    .B2(_05739_),
    .ZN(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05895_ (.A1(_05744_),
    .A2(_05748_),
    .Z(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05896_ (.I(\as2650.r0[2] ),
    .Z(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05897_ (.I(_05750_),
    .Z(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05898_ (.I(_05751_),
    .Z(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05899_ (.I(_05711_),
    .Z(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05900_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_05753_),
    .Z(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _05901_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123[0][2] ),
    .I2(\as2650.r123_2[1][2] ),
    .I3(\as2650.r123_2[0][2] ),
    .S0(_05705_),
    .S1(_05753_),
    .Z(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _05902_ (.A1(_05752_),
    .A2(_05726_),
    .B1(_05754_),
    .B2(_05718_),
    .C1(_05755_),
    .C2(_05706_),
    .ZN(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05903_ (.I(_05756_),
    .Z(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05904_ (.I(\as2650.r0[4] ),
    .Z(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05905_ (.I(_05758_),
    .Z(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05906_ (.I(_05759_),
    .Z(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05907_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_05736_),
    .Z(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _05908_ (.I0(\as2650.r123[1][4] ),
    .I1(\as2650.r123[0][4] ),
    .I2(\as2650.r123_2[1][4] ),
    .I3(\as2650.r123_2[0][4] ),
    .S0(_05683_),
    .S1(_05736_),
    .Z(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _05909_ (.A1(_05760_),
    .A2(_05734_),
    .B1(_05761_),
    .B2(_05719_),
    .C1(_05762_),
    .C2(_05739_),
    .ZN(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05910_ (.I(\as2650.r0[3] ),
    .Z(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05911_ (.I(_05764_),
    .Z(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05912_ (.I(_05765_),
    .Z(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05913_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_05712_),
    .Z(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05914_ (.I0(\as2650.r123[1][3] ),
    .I1(\as2650.r123[0][3] ),
    .I2(\as2650.r123_2[1][3] ),
    .I3(\as2650.r123_2[0][3] ),
    .S0(_05683_),
    .S1(_05712_),
    .Z(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05915_ (.A1(_05766_),
    .A2(_05726_),
    .B1(_05767_),
    .B2(_05718_),
    .C1(_05768_),
    .C2(_05707_),
    .ZN(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05916_ (.I(_05769_),
    .Z(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05917_ (.I(\as2650.alu_op[0] ),
    .Z(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05918_ (.A1(\as2650.alu_op[2] ),
    .A2(\as2650.alu_op[1] ),
    .Z(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05919_ (.A1(\as2650.ins_reg[4] ),
    .A2(_05772_),
    .ZN(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05920_ (.I(\as2650.r0[0] ),
    .Z(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05921_ (.I(_05774_),
    .Z(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05922_ (.I(_05775_),
    .Z(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05923_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(_05711_),
    .Z(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _05924_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123[0][0] ),
    .I2(\as2650.r123_2[1][0] ),
    .I3(\as2650.r123_2[0][0] ),
    .S0(\as2650.ins_reg[0] ),
    .S1(_05711_),
    .Z(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _05925_ (.A1(_05776_),
    .A2(_05725_),
    .B1(_05777_),
    .B2(_05717_),
    .C1(_05778_),
    .C2(_05706_),
    .ZN(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05926_ (.I(\as2650.r0[1] ),
    .Z(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05927_ (.I(_05780_),
    .Z(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05928_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_05753_),
    .Z(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _05929_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123[0][1] ),
    .I2(\as2650.r123_2[1][1] ),
    .I3(\as2650.r123_2[0][1] ),
    .S0(_05705_),
    .S1(_05753_),
    .Z(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _05930_ (.A1(_05781_),
    .A2(_05725_),
    .B1(_05782_),
    .B2(_05717_),
    .C1(_05783_),
    .C2(_05706_),
    .ZN(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05931_ (.A1(_05771_),
    .A2(_05773_),
    .A3(_05779_),
    .A4(_05784_),
    .Z(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05932_ (.A1(_05757_),
    .A2(_05763_),
    .A3(_05770_),
    .A4(_05785_),
    .Z(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05933_ (.A1(\as2650.alu_op[2] ),
    .A2(_05692_),
    .ZN(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05934_ (.A1(\as2650.ins_reg[4] ),
    .A2(\as2650.alu_op[0] ),
    .ZN(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05935_ (.A1(_05787_),
    .A2(_05788_),
    .ZN(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05936_ (.I(_05779_),
    .Z(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05937_ (.A1(_05789_),
    .A2(_05790_),
    .Z(_05791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05938_ (.I(_05784_),
    .Z(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05939_ (.A1(_05757_),
    .A2(_05792_),
    .A3(_05763_),
    .A4(_05769_),
    .Z(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05940_ (.A1(_05741_),
    .A2(_05791_),
    .A3(_05793_),
    .A4(_05749_),
    .ZN(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05941_ (.A1(_05741_),
    .A2(_05749_),
    .A3(_05786_),
    .B(_05794_),
    .ZN(_05795_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05942_ (.A1(_05730_),
    .A2(_05795_),
    .Z(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05943_ (.I(_05749_),
    .Z(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05944_ (.A1(_05791_),
    .A2(_05793_),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05945_ (.A1(_05735_),
    .A2(_05740_),
    .ZN(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05946_ (.I0(_05798_),
    .I1(_05786_),
    .S(_05799_),
    .Z(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05947_ (.A1(_05797_),
    .A2(_05800_),
    .Z(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05948_ (.I(_05799_),
    .Z(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05949_ (.A1(_05798_),
    .A2(_05786_),
    .ZN(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05950_ (.A1(_05802_),
    .A2(_05803_),
    .Z(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05951_ (.A1(_05760_),
    .A2(_05727_),
    .ZN(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05952_ (.A1(_05745_),
    .A2(_05761_),
    .B1(_05762_),
    .B2(_05708_),
    .ZN(_05806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05953_ (.A1(_05805_),
    .A2(_05806_),
    .ZN(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05954_ (.I(_05756_),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05955_ (.I(_05784_),
    .Z(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05956_ (.A1(_05790_),
    .A2(_05757_),
    .A3(_05809_),
    .A4(_05769_),
    .ZN(_05810_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05957_ (.I(_05789_),
    .ZN(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _05958_ (.A1(_05808_),
    .A2(_05770_),
    .A3(_05785_),
    .B1(_05810_),
    .B2(_05811_),
    .ZN(_05812_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05959_ (.A1(_05807_),
    .A2(_05812_),
    .Z(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05960_ (.I(_05752_),
    .Z(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05961_ (.A1(_05814_),
    .A2(_05734_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05962_ (.A1(_05719_),
    .A2(_05754_),
    .B1(_05755_),
    .B2(_05707_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05963_ (.A1(_00420_),
    .A2(_00421_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05964_ (.I(_00422_),
    .Z(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05965_ (.A1(_05789_),
    .A2(_05790_),
    .A3(_05809_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05966_ (.A1(_00424_),
    .A2(_05785_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05967_ (.A1(_00423_),
    .A2(_00425_),
    .Z(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05968_ (.I(_05790_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05969_ (.A1(_05773_),
    .A2(_00427_),
    .Z(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05970_ (.I(_05779_),
    .Z(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05971_ (.I(_00429_),
    .Z(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05972_ (.A1(_05771_),
    .A2(_05773_),
    .A3(_00430_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05973_ (.I(_05792_),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05974_ (.A1(_05791_),
    .A2(_00431_),
    .B(_00432_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05975_ (.I(_05809_),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05976_ (.A1(_05791_),
    .A2(_00434_),
    .A3(_00431_),
    .Z(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05977_ (.A1(_00428_),
    .A2(_00433_),
    .A3(_00435_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05978_ (.I(_05769_),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05979_ (.I0(_00424_),
    .I1(_05785_),
    .S(_00422_),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05980_ (.A1(_00437_),
    .A2(_00438_),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05981_ (.A1(_05813_),
    .A2(_00426_),
    .A3(_00436_),
    .A4(_00439_),
    .Z(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05982_ (.A1(_05796_),
    .A2(_05801_),
    .A3(_05804_),
    .A4(_00440_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05983_ (.A1(_05704_),
    .A2(_05693_),
    .A3(_00441_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05984_ (.A1(_05703_),
    .A2(_00442_),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05985_ (.I(_00443_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05986_ (.I(_00444_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05987_ (.I(_00445_),
    .Z(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05988_ (.I(\as2650.ins_reg[3] ),
    .Z(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05989_ (.I(_00447_),
    .Z(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05990_ (.A1(_00448_),
    .A2(_05700_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05991_ (.I(_00449_),
    .Z(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05992_ (.I(_00450_),
    .Z(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05993_ (.I(_00451_),
    .Z(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05994_ (.I(_05691_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05995_ (.A1(_00453_),
    .A2(_05692_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05996_ (.I(_00447_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05997_ (.A1(_00455_),
    .A2(_05679_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05998_ (.A1(_05720_),
    .A2(_00454_),
    .A3(_00456_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05999_ (.I(_00457_),
    .Z(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06000_ (.I(\as2650.prefixed ),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06001_ (.I(_05771_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06002_ (.I(_05772_),
    .Z(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06003_ (.A1(_00460_),
    .A2(_00461_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06004_ (.I(\as2650.ins_reg[2] ),
    .Z(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06005_ (.A1(_00463_),
    .A2(_00455_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06006_ (.A1(_05700_),
    .A2(_00462_),
    .A3(_00464_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06007_ (.A1(_05728_),
    .A2(_00465_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06008_ (.I(net72),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06009_ (.I(\as2650.cycle[0] ),
    .Z(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06010_ (.A1(_00467_),
    .A2(_00468_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06011_ (.I(_00469_),
    .Z(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06012_ (.A1(_00466_),
    .A2(_00470_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06013_ (.A1(_00459_),
    .A2(_00471_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06014_ (.A1(_00458_),
    .A2(_00472_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06015_ (.I(_00473_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06016_ (.A1(_05678_),
    .A2(_00446_),
    .A3(_00452_),
    .A4(_00474_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06017_ (.I(_05688_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06018_ (.I(_05684_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06019_ (.A1(_00476_),
    .A2(_00477_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06020_ (.A1(_05699_),
    .A2(_00462_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06021_ (.I(_00463_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06022_ (.A1(_00480_),
    .A2(_00447_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06023_ (.A1(_00479_),
    .A2(_00481_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06024_ (.A1(_00478_),
    .A2(_00482_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06025_ (.A1(net72),
    .A2(\as2650.cycle[0] ),
    .Z(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06026_ (.I(_00484_),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06027_ (.A1(_00483_),
    .A2(_00485_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06028_ (.I(\as2650.prefixed ),
    .Z(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06029_ (.A1(_00487_),
    .A2(_00448_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06030_ (.I(_00488_),
    .Z(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06031_ (.A1(_00486_),
    .A2(_00489_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06032_ (.I(_05691_),
    .Z(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06033_ (.I(_00463_),
    .Z(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06034_ (.I(_05788_),
    .Z(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06035_ (.A1(_00492_),
    .A2(_00493_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06036_ (.A1(_00491_),
    .A2(_00494_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06037_ (.I(_00495_),
    .Z(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06038_ (.A1(_05676_),
    .A2(_00496_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06039_ (.I(_00497_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06040_ (.A1(_00490_),
    .A2(_00498_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06041_ (.I(_00453_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06042_ (.A1(_00500_),
    .A2(_00494_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06043_ (.I(_00501_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06044_ (.I(_05699_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06045_ (.A1(_00455_),
    .A2(_00503_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06046_ (.A1(_00487_),
    .A2(_00504_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06047_ (.I(_00505_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06048_ (.A1(_05675_),
    .A2(_00485_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06049_ (.A1(_00506_),
    .A2(_00507_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06050_ (.A1(_00502_),
    .A2(_00508_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06051_ (.I(_05676_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06052_ (.I(_00510_),
    .Z(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06053_ (.I(_00511_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06054_ (.I(_00492_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06055_ (.I(_05720_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06056_ (.I(_00454_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06057_ (.A1(_00514_),
    .A2(_00515_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06058_ (.A1(_00449_),
    .A2(_00516_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06059_ (.A1(_00513_),
    .A2(_00517_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06060_ (.I(_00518_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06061_ (.I(_00519_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06062_ (.I(_00520_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06063_ (.I(_00521_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06064_ (.I(_00456_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06065_ (.A1(_00487_),
    .A2(_00484_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06066_ (.A1(_00523_),
    .A2(_00524_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06067_ (.A1(_00512_),
    .A2(_00522_),
    .A3(_00525_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06068_ (.A1(_00475_),
    .A2(_00499_),
    .A3(_00509_),
    .A4(_00526_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06069_ (.I(net5),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06070_ (.I(_00528_),
    .Z(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06071_ (.I(\as2650.cycle[10] ),
    .Z(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06072_ (.I(net6),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06073_ (.A1(_00530_),
    .A2(\as2650.cycle[2] ),
    .B(_00531_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06074_ (.I(_00532_),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06075_ (.I(_00533_),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06076_ (.I(net6),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06077_ (.I(_00535_),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06078_ (.A1(_00536_),
    .A2(\as2650.cycle[3] ),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06079_ (.I(_00537_),
    .Z(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06080_ (.A1(_00529_),
    .A2(_00534_),
    .A3(_00538_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06081_ (.I(_00531_),
    .Z(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06082_ (.A1(_00540_),
    .A2(\as2650.cycle[11] ),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06083_ (.A1(\as2650.prefixed ),
    .A2(_05699_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06084_ (.A1(_00469_),
    .A2(_00542_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06085_ (.A1(\as2650.cycle[13] ),
    .A2(_00535_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06086_ (.A1(_00543_),
    .A2(_00544_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06087_ (.A1(_00466_),
    .A2(_00545_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06088_ (.A1(_00541_),
    .A2(_00546_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06089_ (.I(_00536_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06090_ (.I(_00548_),
    .Z(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06091_ (.I(\as2650.cycle[1] ),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06092_ (.A1(_00549_),
    .A2(_00550_),
    .Z(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06093_ (.I(_00551_),
    .Z(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06094_ (.A1(_00539_),
    .A2(_00547_),
    .A3(_00552_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06095_ (.A1(_00535_),
    .A2(\as2650.cycle[11] ),
    .Z(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06096_ (.I(_00554_),
    .Z(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06097_ (.I(_00555_),
    .Z(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06098_ (.I(_00466_),
    .Z(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06099_ (.A1(\as2650.cycle[13] ),
    .A2(net6),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06100_ (.I(_00558_),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06101_ (.A1(_00458_),
    .A2(_00557_),
    .A3(_00559_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06102_ (.I(\as2650.cycle[5] ),
    .Z(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06103_ (.A1(_00531_),
    .A2(_00561_),
    .Z(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06104_ (.A1(_00525_),
    .A2(_00562_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06105_ (.I(\as2650.cycle[4] ),
    .Z(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06106_ (.A1(_00536_),
    .A2(_00564_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06107_ (.A1(_00563_),
    .A2(_00565_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06108_ (.A1(_00560_),
    .A2(_00566_),
    .Z(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06109_ (.I(net7),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06110_ (.A1(_00568_),
    .A2(\as2650.last_intr ),
    .A3(net75),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06111_ (.A1(_00467_),
    .A2(_00569_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06112_ (.I(_00570_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06113_ (.A1(_00485_),
    .A2(_00571_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06114_ (.A1(_00549_),
    .A2(\as2650.cycle[7] ),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06115_ (.I(_00524_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06116_ (.A1(_00535_),
    .A2(_00561_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06117_ (.I(_00575_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06118_ (.A1(_00523_),
    .A2(_00574_),
    .A3(_00576_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06119_ (.A1(_00480_),
    .A2(_00457_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06120_ (.A1(_00578_),
    .A2(_00559_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06121_ (.I(_00579_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06122_ (.A1(_00540_),
    .A2(\as2650.cycle[12] ),
    .Z(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06123_ (.A1(_00577_),
    .A2(_00580_),
    .A3(_00581_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06124_ (.A1(_00573_),
    .A2(_00582_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06125_ (.A1(_00556_),
    .A2(_00567_),
    .B(_00572_),
    .C(_00583_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06126_ (.I(_00544_),
    .Z(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06127_ (.I(_00585_),
    .Z(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06128_ (.A1(_00463_),
    .A2(_05679_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06129_ (.I(_00587_),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06130_ (.I(_05771_),
    .Z(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06131_ (.I(_00589_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06132_ (.A1(_00453_),
    .A2(_05692_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06133_ (.I(_00591_),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06134_ (.A1(_00590_),
    .A2(_00592_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06135_ (.A1(_00588_),
    .A2(_00593_),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06136_ (.A1(_00589_),
    .A2(_05787_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06137_ (.A1(_00595_),
    .A2(_00587_),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06138_ (.A1(_00594_),
    .A2(_00596_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06139_ (.I(_00597_),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06140_ (.A1(_00496_),
    .A2(_00598_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06141_ (.A1(_00508_),
    .A2(_00599_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06142_ (.I(_00480_),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06143_ (.A1(_00601_),
    .A2(_05702_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06144_ (.A1(_00494_),
    .A2(_00602_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06145_ (.A1(_00600_),
    .A2(_00603_),
    .B(_00509_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06146_ (.I(_00459_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06147_ (.I(_00605_),
    .Z(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06148_ (.A1(_00601_),
    .A2(_00517_),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06149_ (.I(_00607_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06150_ (.A1(_00489_),
    .A2(_00594_),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06151_ (.A1(_00606_),
    .A2(_00608_),
    .A3(_00585_),
    .B(_00609_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06152_ (.I(_00595_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06153_ (.A1(_00611_),
    .A2(_00588_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06154_ (.I(_00612_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06155_ (.A1(_00492_),
    .A2(_00503_),
    .A3(_05701_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06156_ (.I(_00614_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06157_ (.I(_00615_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06158_ (.A1(_00613_),
    .A2(_00616_),
    .B(_00508_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06159_ (.A1(_00507_),
    .A2(_00610_),
    .B(_00617_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06160_ (.A1(_00586_),
    .A2(_00604_),
    .B(_00618_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06161_ (.A1(_00529_),
    .A2(_00584_),
    .B(_00619_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06162_ (.I(_00620_),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06163_ (.I(\as2650.cycle[13] ),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06164_ (.I(_00622_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06165_ (.A1(_00553_),
    .A2(_00621_),
    .B(_00623_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06166_ (.I(_00547_),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06167_ (.I(net3),
    .Z(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06168_ (.I(_00626_),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06169_ (.I(_00627_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06170_ (.I(_00628_),
    .Z(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06171_ (.I(_00629_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06172_ (.A1(_00536_),
    .A2(\as2650.cycle[1] ),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06173_ (.I(_00631_),
    .Z(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06174_ (.I(_00632_),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06175_ (.A1(\as2650.cycle[9] ),
    .A2(_00632_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06176_ (.A1(_00511_),
    .A2(_00630_),
    .A3(_00633_),
    .B1(_00634_),
    .B2(_00539_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06177_ (.I(_00635_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06178_ (.I(\as2650.addr_buff[7] ),
    .Z(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06179_ (.I(_00637_),
    .Z(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06180_ (.I(_00638_),
    .Z(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06181_ (.I(_00510_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06182_ (.A1(_00540_),
    .A2(_00530_),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06183_ (.A1(_00641_),
    .A2(_00537_),
    .A3(_00631_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06184_ (.A1(_00639_),
    .A2(_00640_),
    .A3(_00547_),
    .A4(_00642_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06185_ (.A1(_00625_),
    .A2(_00636_),
    .B(_00643_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06186_ (.I(_05669_),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06187_ (.A1(_00645_),
    .A2(_05675_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06188_ (.I(_00542_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06189_ (.I(_00494_),
    .Z(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06190_ (.A1(_00588_),
    .A2(_00593_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06191_ (.A1(_00649_),
    .A2(_00612_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06192_ (.I(_05728_),
    .Z(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06193_ (.A1(_00460_),
    .A2(_00454_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06194_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06195_ (.I(_00653_),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06196_ (.I(_00654_),
    .Z(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06197_ (.I(_00655_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06198_ (.A1(_05680_),
    .A2(_00652_),
    .A3(_00656_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06199_ (.A1(_00651_),
    .A2(_00657_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06200_ (.A1(_00486_),
    .A2(_00505_),
    .A3(_00614_),
    .A4(_00658_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06201_ (.A1(_00648_),
    .A2(_00650_),
    .A3(_00659_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06202_ (.A1(_00647_),
    .A2(_00660_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06203_ (.I(_00486_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06204_ (.I(_00589_),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06205_ (.A1(\as2650.ins_reg[2] ),
    .A2(_00447_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06206_ (.I(_00664_),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06207_ (.I(_00665_),
    .Z(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06208_ (.I(_00666_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06209_ (.A1(_00651_),
    .A2(_00667_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06210_ (.A1(_05704_),
    .A2(_00663_),
    .A3(_05694_),
    .A4(_00668_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06211_ (.A1(_00500_),
    .A2(_00669_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06212_ (.A1(_00662_),
    .A2(_00670_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06213_ (.I(_00608_),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06214_ (.I(_00672_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06215_ (.A1(_00464_),
    .A2(_00661_),
    .A3(_00671_),
    .B1(_00673_),
    .B2(_00525_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06216_ (.A1(_00462_),
    .A2(_00644_),
    .B1(_00646_),
    .B2(_00674_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06217_ (.A1(_05674_),
    .A2(_00527_),
    .B(_00624_),
    .C(_00675_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06218_ (.A1(_00472_),
    .A2(_00673_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06219_ (.I(_00529_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06220_ (.I(_00677_),
    .Z(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06221_ (.I(_00523_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06222_ (.I(_00679_),
    .Z(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06223_ (.I(_00562_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06224_ (.A1(_00638_),
    .A2(_00681_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06225_ (.I(_00682_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06226_ (.A1(_00678_),
    .A2(_00680_),
    .A3(_00683_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06227_ (.A1(_00448_),
    .A2(_05680_),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06228_ (.A1(_00524_),
    .A2(_00685_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06229_ (.I(_00562_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06230_ (.I(_00687_),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06231_ (.I(_00688_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06232_ (.A1(_00498_),
    .A2(_00686_),
    .A3(_00689_),
    .B(_00620_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06233_ (.A1(_00553_),
    .A2(_00690_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06234_ (.I(_00691_),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06235_ (.A1(\as2650.cycle[12] ),
    .A2(_00692_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06236_ (.A1(_00676_),
    .A2(_00580_),
    .A3(_00684_),
    .B(_00693_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06237_ (.I(\as2650.cycle[4] ),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06238_ (.I(_00510_),
    .Z(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06239_ (.I(_00695_),
    .Z(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06240_ (.I(_00696_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06241_ (.I(_00576_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06242_ (.I(_00698_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06243_ (.A1(_00520_),
    .A2(_00699_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06244_ (.A1(_00492_),
    .A2(_00457_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06245_ (.I(_00701_),
    .Z(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06246_ (.I(_00544_),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06247_ (.A1(_00702_),
    .A2(_00703_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06248_ (.A1(_00679_),
    .A2(_00574_),
    .A3(_00704_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06249_ (.A1(_00700_),
    .A2(_00705_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06250_ (.I(_00549_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06251_ (.A1(_00482_),
    .A2(_00545_),
    .B1(_00706_),
    .B2(_00707_),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06252_ (.I(\as2650.cycle[11] ),
    .Z(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06253_ (.A1(_00709_),
    .A2(_00692_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06254_ (.A1(_00694_),
    .A2(_00697_),
    .A3(_00708_),
    .B(_00710_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06255_ (.I(_00640_),
    .Z(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06256_ (.I(_00711_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06257_ (.I(\as2650.cycle[3] ),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06258_ (.A1(_00548_),
    .A2(_00713_),
    .Z(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06259_ (.A1(_00714_),
    .A2(_00632_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06260_ (.A1(_00530_),
    .A2(_00692_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06261_ (.A1(_00712_),
    .A2(_00625_),
    .A3(_00715_),
    .B(_00716_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06262_ (.I(_00551_),
    .Z(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06263_ (.I(_00714_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06264_ (.I(_00718_),
    .Z(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06265_ (.I(\as2650.cycle[2] ),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06266_ (.A1(_00531_),
    .A2(\as2650.cycle[10] ),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06267_ (.I(_00721_),
    .Z(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06268_ (.A1(_00549_),
    .A2(_00720_),
    .A3(_00722_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06269_ (.A1(_00711_),
    .A2(_00719_),
    .A3(_00723_),
    .Z(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06270_ (.I(\as2650.cycle[9] ),
    .Z(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06271_ (.A1(_00725_),
    .A2(_00690_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06272_ (.A1(_00625_),
    .A2(_00717_),
    .A3(_00724_),
    .B(_00726_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06273_ (.I(_05678_),
    .Z(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06274_ (.I(_00727_),
    .Z(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06275_ (.I(_00470_),
    .Z(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06276_ (.I(_00729_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06277_ (.I(_00730_),
    .Z(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06278_ (.I(_00731_),
    .Z(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06279_ (.A1(_00707_),
    .A2(_00732_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06280_ (.I(\as2650.cycle[8] ),
    .Z(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06281_ (.I(_00734_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06282_ (.I(_00735_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06283_ (.I(_00736_),
    .Z(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06284_ (.A1(_00468_),
    .A2(_00570_),
    .B1(_00733_),
    .B2(_00737_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06285_ (.A1(_00728_),
    .A2(_00738_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06286_ (.I(_00711_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06287_ (.A1(_00518_),
    .A2(_00681_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06288_ (.A1(_00581_),
    .A2(_00740_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06289_ (.A1(\as2650.cycle[7] ),
    .A2(_00691_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06290_ (.A1(_00739_),
    .A2(_00705_),
    .A3(_00741_),
    .B(_00742_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06291_ (.I(\as2650.cycle[6] ),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06292_ (.A1(_00743_),
    .A2(_00528_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06293_ (.I(_00744_),
    .Z(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06294_ (.I(\as2650.cycle[8] ),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06295_ (.I(_00746_),
    .Z(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06296_ (.I(_00485_),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06297_ (.I(_00748_),
    .Z(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06298_ (.A1(_00747_),
    .A2(_05678_),
    .A3(_00749_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06299_ (.I(_00750_),
    .Z(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06300_ (.A1(_00707_),
    .A2(_00751_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06301_ (.A1(_00572_),
    .A2(_00745_),
    .B(_00752_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06302_ (.A1(_00662_),
    .A2(_00608_),
    .A3(_00585_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06303_ (.I(_00606_),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06304_ (.I(_00754_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06305_ (.I(_00755_),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06306_ (.I(_00756_),
    .Z(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06307_ (.I(_00685_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06308_ (.I(_00758_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06309_ (.I(_00759_),
    .Z(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06310_ (.A1(_00757_),
    .A2(_00696_),
    .A3(_00588_),
    .A4(_00760_),
    .Z(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06311_ (.I(_00671_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06312_ (.I(_00479_),
    .Z(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06313_ (.I(_00656_),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06314_ (.I(_00764_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06315_ (.I(_05701_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06316_ (.A1(_05704_),
    .A2(_00590_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06317_ (.A1(_00766_),
    .A2(_00767_),
    .Z(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06318_ (.I(_00768_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06319_ (.A1(_00647_),
    .A2(_00646_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06320_ (.A1(_00763_),
    .A2(_00765_),
    .A3(_00769_),
    .A4(_00770_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06321_ (.I(\as2650.cycle[5] ),
    .Z(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06322_ (.I(_00772_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06323_ (.I(_00773_),
    .Z(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06324_ (.I(_00774_),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _06325_ (.A1(_00623_),
    .A2(_00499_),
    .B1(_00762_),
    .B2(_00771_),
    .C1(_00690_),
    .C2(_00775_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06326_ (.A1(_00753_),
    .A2(_00761_),
    .B(_00776_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06327_ (.A1(_00564_),
    .A2(_00690_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06328_ (.I(_00513_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06329_ (.I(_00778_),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06330_ (.I(_00779_),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06331_ (.I(_00780_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06332_ (.I(_00458_),
    .Z(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06333_ (.I(_00782_),
    .Z(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06334_ (.I(_00559_),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06335_ (.I(_00784_),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06336_ (.I(_00785_),
    .Z(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06337_ (.I(_00786_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06338_ (.A1(_00781_),
    .A2(_00783_),
    .A3(_00787_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06339_ (.I(_00451_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06340_ (.A1(_00781_),
    .A2(_00789_),
    .A3(_00474_),
    .A4(_00787_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06341_ (.A1(_00574_),
    .A2(_00788_),
    .B(_00790_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06342_ (.I(net3),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06343_ (.I(_00792_),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06344_ (.I(_00793_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06345_ (.I(_00794_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _06346_ (.A1(_00474_),
    .A2(_00586_),
    .A3(_00684_),
    .B1(_00791_),
    .B2(_00512_),
    .B3(_00795_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06347_ (.A1(_00611_),
    .A2(_00644_),
    .B(_00796_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06348_ (.A1(_00777_),
    .A2(_00797_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06349_ (.I(_00448_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06350_ (.I(_00798_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06351_ (.I(_00799_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06352_ (.I(_00800_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06353_ (.A1(_00781_),
    .A2(_00801_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06354_ (.A1(_00713_),
    .A2(_00691_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06355_ (.A1(_00671_),
    .A2(_00802_),
    .A3(_00770_),
    .B(_00803_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06356_ (.I(_00601_),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06357_ (.I(_00804_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06358_ (.A1(_00805_),
    .A2(_00801_),
    .A3(_00646_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06359_ (.A1(_00550_),
    .A2(_00692_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06360_ (.A1(_00543_),
    .A2(_00806_),
    .B(_00807_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06361_ (.I(_00627_),
    .Z(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06362_ (.I(_00808_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06363_ (.I(_00809_),
    .Z(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06364_ (.I(_00810_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06365_ (.A1(_00550_),
    .A2(_00713_),
    .A3(_00721_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06366_ (.A1(_00811_),
    .A2(_00717_),
    .B1(_00812_),
    .B2(_00639_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06367_ (.A1(_00720_),
    .A2(_00691_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06368_ (.A1(_00739_),
    .A2(_00625_),
    .A3(_00813_),
    .B(_00814_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06369_ (.A1(_00607_),
    .A2(_00559_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06370_ (.I(_00815_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06371_ (.A1(\as2650.addr_buff[7] ),
    .A2(_00575_),
    .Z(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06372_ (.I(_00817_),
    .Z(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06373_ (.A1(_00512_),
    .A2(_00816_),
    .A3(_00818_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06374_ (.A1(_00474_),
    .A2(_00745_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06375_ (.A1(_00472_),
    .A2(_00819_),
    .B1(_00820_),
    .B2(_00446_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06376_ (.I(_00731_),
    .Z(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06377_ (.I(_00755_),
    .Z(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06378_ (.I(_00823_),
    .Z(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06379_ (.I(_00491_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06380_ (.I(_00477_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06381_ (.I(_05693_),
    .Z(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06382_ (.I(_00653_),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06383_ (.I(_00828_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06384_ (.I(_00829_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06385_ (.A1(_05696_),
    .A2(_00830_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06386_ (.A1(_00826_),
    .A2(_00827_),
    .A3(_00767_),
    .A4(_00831_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06387_ (.A1(_00825_),
    .A2(_00832_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06388_ (.I(_00658_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06389_ (.I(_00834_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06390_ (.A1(_00511_),
    .A2(_00835_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06391_ (.I(_05685_),
    .Z(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06392_ (.A1(_00476_),
    .A2(_00837_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06393_ (.A1(_00590_),
    .A2(_05695_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06394_ (.A1(_00503_),
    .A2(_00839_),
    .A3(_00667_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06395_ (.A1(_00838_),
    .A2(_00840_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06396_ (.I(_00841_),
    .Z(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06397_ (.I(_00837_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06398_ (.A1(_00590_),
    .A2(_05702_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06399_ (.I(_00844_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06400_ (.A1(_00831_),
    .A2(_00845_),
    .ZN(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06401_ (.A1(_00843_),
    .A2(_00846_),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06402_ (.A1(_00842_),
    .A2(_00847_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06403_ (.I(_00667_),
    .Z(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06404_ (.A1(_00514_),
    .A2(_00849_),
    .A3(_00845_),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06405_ (.A1(_00476_),
    .A2(_00843_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06406_ (.A1(_00851_),
    .A2(_00657_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06407_ (.I(_00852_),
    .Z(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06408_ (.A1(_00848_),
    .A2(_00850_),
    .A3(_00853_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06409_ (.A1(_05701_),
    .A2(_00767_),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06410_ (.A1(_00511_),
    .A2(_00765_),
    .A3(_00855_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06411_ (.A1(_00833_),
    .A2(_00836_),
    .A3(_00854_),
    .A4(_00856_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06412_ (.A1(_00824_),
    .A2(_00857_),
    .B(_00609_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06413_ (.A1(_00831_),
    .A2(_00844_),
    .Z(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06414_ (.A1(_00843_),
    .A2(_00859_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06415_ (.I(_00860_),
    .Z(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06416_ (.I(\as2650.prefixed ),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06417_ (.I(_00862_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06418_ (.I(_00863_),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06419_ (.I(_00864_),
    .Z(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06420_ (.I(_00651_),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06421_ (.A1(_00866_),
    .A2(_00763_),
    .A3(_00849_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06422_ (.A1(_00865_),
    .A2(_00677_),
    .A3(_00763_),
    .A4(_00867_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06423_ (.A1(_00765_),
    .A2(_00671_),
    .A3(_00768_),
    .A4(_00868_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06424_ (.A1(_00505_),
    .A2(_00834_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06425_ (.I(_00666_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06426_ (.I(_00871_),
    .Z(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06427_ (.A1(_00851_),
    .A2(_00872_),
    .A3(_00845_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06428_ (.I(_00873_),
    .Z(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06429_ (.A1(_00471_),
    .A2(_00870_),
    .A3(_00874_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06430_ (.A1(_00543_),
    .A2(_00867_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06431_ (.A1(_00617_),
    .A2(_00869_),
    .A3(_00875_),
    .A4(_00876_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06432_ (.I(_05704_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06433_ (.I(_00878_),
    .Z(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06434_ (.I(_00879_),
    .Z(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06435_ (.I(_00880_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06436_ (.I(_00881_),
    .Z(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06437_ (.I(_00849_),
    .Z(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06438_ (.I(_00663_),
    .Z(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06439_ (.I(_00884_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06440_ (.I(_00885_),
    .Z(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06441_ (.A1(_00886_),
    .A2(_00516_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06442_ (.A1(_00882_),
    .A2(_00883_),
    .A3(_00660_),
    .A4(_00887_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06443_ (.A1(_00659_),
    .A2(_00861_),
    .B(_00877_),
    .C(_00888_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06444_ (.A1(_00822_),
    .A2(_00858_),
    .B(_00889_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06445_ (.A1(_00557_),
    .A2(_00545_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06446_ (.A1(_00891_),
    .A2(_00567_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06447_ (.I(_00576_),
    .Z(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06448_ (.I(_00893_),
    .Z(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06449_ (.I(_00894_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06450_ (.I(_00895_),
    .Z(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06451_ (.A1(_00686_),
    .A2(_00896_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06452_ (.A1(_00589_),
    .A2(_00587_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06453_ (.A1(_00500_),
    .A2(_00898_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06454_ (.A1(_00468_),
    .A2(_00571_),
    .B1(_00897_),
    .B2(_00899_),
    .C(_05678_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06455_ (.A1(_00862_),
    .A2(_00557_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06456_ (.A1(_00720_),
    .A2(_00725_),
    .A3(\as2650.cycle[12] ),
    .A4(\as2650.cycle[7] ),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06457_ (.A1(_00468_),
    .A2(_00550_),
    .A3(_00713_),
    .A4(_00530_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06458_ (.A1(\as2650.cycle[4] ),
    .A2(_00561_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06459_ (.A1(_00645_),
    .A2(_00904_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06460_ (.I(_00905_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06461_ (.A1(_00623_),
    .A2(_00709_),
    .A3(_00903_),
    .A4(_00906_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06462_ (.A1(_00902_),
    .A2(_00907_),
    .B(_05677_),
    .C(_00749_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06463_ (.A1(_00509_),
    .A2(_00586_),
    .B1(_00901_),
    .B2(_00908_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06464_ (.A1(_00577_),
    .A2(_00573_),
    .A3(_00580_),
    .A4(_00581_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06465_ (.I(_00466_),
    .Z(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06466_ (.A1(_00911_),
    .A2(_00501_),
    .A3(_00703_),
    .A4(_00615_),
    .ZN(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06467_ (.A1(_00694_),
    .A2(_00510_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06468_ (.I(_00774_),
    .Z(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06469_ (.A1(_00465_),
    .A2(_00913_),
    .B(_00914_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06470_ (.A1(_00508_),
    .A2(_00599_),
    .A3(_00912_),
    .B1(_00915_),
    .B2(_00891_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06471_ (.A1(_00910_),
    .A2(_00916_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06472_ (.A1(_00900_),
    .A2(_00909_),
    .A3(_00917_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06473_ (.A1(_00512_),
    .A2(_00811_),
    .A3(_00791_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06474_ (.A1(_00556_),
    .A2(_00892_),
    .B(_00918_),
    .C(_00919_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06475_ (.A1(_00452_),
    .A2(_00821_),
    .B1(_00890_),
    .B2(_05674_),
    .C(_00920_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06476_ (.I(net28),
    .ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06477_ (.I(_00851_),
    .Z(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06478_ (.A1(_00491_),
    .A2(_00898_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06479_ (.I(_00922_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06480_ (.A1(_05714_),
    .A2(_05728_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06481_ (.A1(\as2650.cycle[8] ),
    .A2(_00484_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06482_ (.A1(_00529_),
    .A2(_00925_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06483_ (.A1(_00558_),
    .A2(_00926_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06484_ (.I(_00743_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06485_ (.I(_00455_),
    .Z(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06486_ (.A1(_00862_),
    .A2(_00929_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06487_ (.A1(_00928_),
    .A2(_00930_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06488_ (.A1(_00923_),
    .A2(_00924_),
    .A3(_00927_),
    .A4(_00931_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06489_ (.I(_00932_),
    .Z(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06490_ (.I(_00933_),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06491_ (.A1(_00479_),
    .A2(_00872_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06492_ (.A1(_00746_),
    .A2(_00469_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06493_ (.I(_00936_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06494_ (.A1(_00459_),
    .A2(_00937_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06495_ (.A1(_00646_),
    .A2(_00938_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06496_ (.I(_05714_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06497_ (.I(_00478_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06498_ (.A1(_00940_),
    .A2(_00941_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06499_ (.A1(_00935_),
    .A2(_00939_),
    .A3(_00942_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06500_ (.I(_00943_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06501_ (.A1(_00744_),
    .A2(_00937_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06502_ (.I(_00924_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06503_ (.A1(_00945_),
    .A2(_00946_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06504_ (.I(_00487_),
    .Z(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06505_ (.A1(_00948_),
    .A2(_00449_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06506_ (.I(_00949_),
    .Z(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06507_ (.I(_00650_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06508_ (.I(_00489_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06509_ (.A1(_00827_),
    .A2(_00950_),
    .B1(_00951_),
    .B2(_00952_),
    .ZN(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06510_ (.A1(_00947_),
    .A2(_00953_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06511_ (.I(_05714_),
    .Z(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06512_ (.A1(_00645_),
    .A2(_00558_),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06513_ (.I(_00956_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06514_ (.A1(_00663_),
    .A2(_00461_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06515_ (.A1(_00772_),
    .A2(_00958_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06516_ (.I(\as2650.idx_ctrl[1] ),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06517_ (.A1(_00960_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06518_ (.A1(_00478_),
    .A2(_00961_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06519_ (.A1(_00872_),
    .A2(_00959_),
    .A3(_00962_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06520_ (.A1(_00862_),
    .A2(_05680_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06521_ (.A1(_00964_),
    .A2(_00926_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06522_ (.I(_00965_),
    .Z(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06523_ (.A1(_00963_),
    .A2(_00966_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06524_ (.A1(_00955_),
    .A2(_00957_),
    .A3(_00967_),
    .ZN(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06525_ (.A1(_00944_),
    .A2(_00954_),
    .A3(_00968_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06526_ (.I(_00946_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06527_ (.I(_00561_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06528_ (.A1(_00694_),
    .A2(_00971_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06529_ (.I(_00972_),
    .Z(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06530_ (.A1(net5),
    .A2(_00936_),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06531_ (.A1(_00542_),
    .A2(_00974_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06532_ (.I(\as2650.addr_buff[6] ),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06533_ (.I(\as2650.addr_buff[5] ),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06534_ (.I(_00977_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06535_ (.A1(_00976_),
    .A2(_00978_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06536_ (.A1(\as2650.addr_buff[7] ),
    .A2(_00979_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06537_ (.A1(_00973_),
    .A2(_00975_),
    .A3(_00980_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06538_ (.I(_00956_),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06539_ (.A1(_00709_),
    .A2(_00642_),
    .A3(_00982_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06540_ (.A1(_00970_),
    .A2(_00981_),
    .A3(_00983_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06541_ (.I(\as2650.cycle[9] ),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06542_ (.A1(_00537_),
    .A2(_00631_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06543_ (.A1(_00985_),
    .A2(_00554_),
    .A3(_00986_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06544_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(\as2650.idx_ctrl[0] ),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06545_ (.I(_00988_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06546_ (.I(_00989_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06547_ (.I(_00990_),
    .Z(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06548_ (.I(_00743_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06549_ (.A1(_00992_),
    .A2(_00544_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06550_ (.A1(_00532_),
    .A2(_00991_),
    .A3(_00993_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06551_ (.A1(_00972_),
    .A2(_00975_),
    .A3(_00994_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06552_ (.A1(_00970_),
    .A2(_00987_),
    .A3(_00995_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06553_ (.A1(_00934_),
    .A2(_00969_),
    .A3(_00984_),
    .A4(_00996_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06554_ (.A1(_00921_),
    .A2(_00997_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06555_ (.I(_00998_),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06556_ (.I(_00968_),
    .Z(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06557_ (.I(_00946_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06558_ (.I(_00961_),
    .Z(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06559_ (.A1(_00714_),
    .A2(_00555_),
    .A3(_00973_),
    .A4(_01002_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06560_ (.A1(_00540_),
    .A2(_00720_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06561_ (.A1(_00722_),
    .A2(_01004_),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06562_ (.A1(_01005_),
    .A2(_00634_),
    .A3(_00957_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06563_ (.A1(_01001_),
    .A2(_00966_),
    .A3(_01003_),
    .A4(_01006_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06564_ (.I(_00960_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06565_ (.I(\as2650.idx_ctrl[0] ),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06566_ (.A1(_01008_),
    .A2(_01009_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06567_ (.I(_01010_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06568_ (.A1(_00427_),
    .A2(_01011_),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06569_ (.A1(_01001_),
    .A2(_00981_),
    .A3(_00983_),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06570_ (.I(_01013_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06571_ (.I(_00429_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06572_ (.I(\as2650.addr_buff[6] ),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06573_ (.A1(_01016_),
    .A2(_00977_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06574_ (.A1(_01015_),
    .A2(_01017_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06575_ (.I(_01018_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06576_ (.I(_05776_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06577_ (.I(_01020_),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06578_ (.I(_01021_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06579_ (.A1(_01022_),
    .A2(_00944_),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06580_ (.I(_00937_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06581_ (.A1(_00745_),
    .A2(_01024_),
    .A3(_00942_),
    .ZN(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06582_ (.A1(_00930_),
    .A2(_00612_),
    .ZN(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06583_ (.A1(_01025_),
    .A2(_01026_),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06584_ (.I(net50),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06585_ (.I(_05730_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06586_ (.I(net78),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06587_ (.A1(net50),
    .A2(_01030_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06588_ (.A1(_01028_),
    .A2(_01029_),
    .B(_01031_),
    .ZN(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06589_ (.A1(_01027_),
    .A2(_01032_),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06590_ (.I(_00432_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06591_ (.A1(_00609_),
    .A2(_00947_),
    .ZN(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06592_ (.I(_01035_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06593_ (.I(_00596_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06594_ (.A1(_00489_),
    .A2(_01037_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06595_ (.A1(_00947_),
    .A2(_01038_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06596_ (.I(_01039_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06597_ (.I(net8),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06598_ (.I(_01041_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06599_ (.I(_01042_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06600_ (.A1(_00923_),
    .A2(_00946_),
    .A3(_00927_),
    .A4(_00931_),
    .Z(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06601_ (.I(_01044_),
    .Z(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06602_ (.I(_01035_),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06603_ (.A1(_00428_),
    .A2(_01044_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06604_ (.A1(_01043_),
    .A2(_01045_),
    .B(_01046_),
    .C(_01047_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06605_ (.A1(_01034_),
    .A2(_01036_),
    .B(_01040_),
    .C(_01048_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06606_ (.A1(_00935_),
    .A2(_00939_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06607_ (.A1(_01001_),
    .A2(_01050_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06608_ (.I(_01051_),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06609_ (.A1(_01033_),
    .A2(_01049_),
    .B(_01052_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06610_ (.A1(_01013_),
    .A2(_01023_),
    .A3(_01053_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06611_ (.A1(_00970_),
    .A2(_00987_),
    .A3(_00995_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06612_ (.A1(_01014_),
    .A2(_01019_),
    .B(_01054_),
    .C(_01055_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06613_ (.A1(_01007_),
    .A2(_01012_),
    .B(_01056_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06614_ (.I(_00652_),
    .Z(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06615_ (.I(_01058_),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06616_ (.A1(net50),
    .A2(net78),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06617_ (.I(\as2650.holding_reg[0] ),
    .Z(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06618_ (.A1(_01015_),
    .A2(_00665_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06619_ (.A1(_05720_),
    .A2(_05777_),
    .B1(_05778_),
    .B2(_05708_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06620_ (.I(_00988_),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06621_ (.I(_05734_),
    .Z(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06622_ (.A1(_01065_),
    .A2(_00989_),
    .B(_01021_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06623_ (.I(_00653_),
    .Z(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06624_ (.A1(_01063_),
    .A2(_01064_),
    .B(_01066_),
    .C(_01067_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06625_ (.A1(_01061_),
    .A2(_01062_),
    .A3(_01068_),
    .Z(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06626_ (.A1(_01061_),
    .A2(_01067_),
    .Z(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06627_ (.A1(\as2650.holding_reg[0] ),
    .A2(_00654_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06628_ (.A1(_01015_),
    .A2(_00828_),
    .B(_01071_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06629_ (.A1(_01068_),
    .A2(_01070_),
    .B(_01072_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06630_ (.A1(_01069_),
    .A2(_01073_),
    .ZN(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06631_ (.A1(_01060_),
    .A2(_01074_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06632_ (.A1(_01059_),
    .A2(_01075_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06633_ (.A1(_00884_),
    .A2(_00515_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06634_ (.A1(_01031_),
    .A2(_01074_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06635_ (.A1(_01077_),
    .A2(_01078_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06636_ (.I(_00663_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06637_ (.A1(_01080_),
    .A2(_00766_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06638_ (.I(_01081_),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06639_ (.A1(_01061_),
    .A2(_01062_),
    .A3(_01068_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06640_ (.I(_01073_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06641_ (.A1(_01083_),
    .A2(_01084_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06642_ (.I(_00593_),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06643_ (.A1(_00460_),
    .A2(_00591_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06644_ (.I(_01087_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06645_ (.A1(_01086_),
    .A2(_01069_),
    .B1(_01084_),
    .B2(_01088_),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06646_ (.I(_05695_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06647_ (.I(_05694_),
    .Z(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06648_ (.A1(_01080_),
    .A2(_01091_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06649_ (.A1(_01090_),
    .A2(_00592_),
    .A3(_01092_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06650_ (.I(_01093_),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06651_ (.A1(_01082_),
    .A2(_01085_),
    .B(_01089_),
    .C(_01094_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06652_ (.I(_01093_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _06653_ (.A1(_01076_),
    .A2(_01079_),
    .A3(_01095_),
    .B1(_01072_),
    .B2(_01096_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06654_ (.A1(_01000_),
    .A2(_01097_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06655_ (.A1(_01000_),
    .A2(_01057_),
    .B(_01098_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06656_ (.I(_01022_),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06657_ (.I(_01100_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06658_ (.I(_01101_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06659_ (.I(_00955_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06660_ (.I(_00939_),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06661_ (.A1(_01103_),
    .A2(_00835_),
    .A3(_01104_),
    .ZN(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06662_ (.I(_01105_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06663_ (.I(_01106_),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06664_ (.I0(\as2650.r123[0][0] ),
    .I1(\as2650.r123_2[0][0] ),
    .S(_05710_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06665_ (.I(_01108_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06666_ (.I(_01109_),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06667_ (.I(_01110_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06668_ (.I(_01111_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06669_ (.A1(_01102_),
    .A2(_01107_),
    .A3(_01112_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06670_ (.I(_00998_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06671_ (.A1(_00695_),
    .A2(_01106_),
    .A3(_01114_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06672_ (.I(_01115_),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06673_ (.A1(\as2650.r123[1][0] ),
    .A2(_01116_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06674_ (.A1(_00999_),
    .A2(_01099_),
    .B(_01113_),
    .C(_01117_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06675_ (.A1(_00429_),
    .A2(_05809_),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06676_ (.I(_01118_),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06677_ (.I(_00429_),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06678_ (.I(_01009_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06679_ (.A1(_00960_),
    .A2(_01121_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06680_ (.A1(_00960_),
    .A2(_01121_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06681_ (.A1(_01120_),
    .A2(_01122_),
    .B(_01123_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06682_ (.A1(_01119_),
    .A2(_01124_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06683_ (.A1(_01119_),
    .A2(_01124_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06684_ (.A1(_01125_),
    .A2(_01126_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06685_ (.A1(_00637_),
    .A2(_00979_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06686_ (.A1(_00904_),
    .A2(_00965_),
    .A3(_01128_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06687_ (.I(_00993_),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06688_ (.A1(_00541_),
    .A2(_00812_),
    .A3(_01130_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06689_ (.A1(_00942_),
    .A2(_01129_),
    .A3(_01131_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06690_ (.I(_01132_),
    .Z(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06691_ (.I(_05781_),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06692_ (.I(_01134_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06693_ (.I(_01135_),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06694_ (.I(_00943_),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06695_ (.I(_01120_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06696_ (.I(_01138_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06697_ (.I(_01039_),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06698_ (.I(net9),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06699_ (.I(_01141_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06700_ (.A1(_00930_),
    .A2(_00649_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06701_ (.A1(_01143_),
    .A2(_01025_),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06702_ (.I(_01144_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06703_ (.A1(_00433_),
    .A2(_00435_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06704_ (.I(_00932_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06705_ (.A1(_01146_),
    .A2(_01147_),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06706_ (.A1(_01142_),
    .A2(_00934_),
    .B(_01145_),
    .C(_01148_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06707_ (.I(_00423_),
    .Z(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06708_ (.A1(_01150_),
    .A2(_01046_),
    .B(_01040_),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06709_ (.A1(_01139_),
    .A2(_01140_),
    .B1(_01149_),
    .B2(_01151_),
    .C(_00943_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06710_ (.A1(_01136_),
    .A2(_01137_),
    .B(_01152_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06711_ (.I(_01132_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06712_ (.I(\as2650.addr_buff[5] ),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06713_ (.A1(_00976_),
    .A2(_01155_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06714_ (.A1(_00976_),
    .A2(_01155_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06715_ (.A1(_01120_),
    .A2(_01156_),
    .B(_01157_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06716_ (.A1(_01119_),
    .A2(_01158_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06717_ (.A1(_01119_),
    .A2(_01158_),
    .ZN(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06718_ (.A1(_01159_),
    .A2(_01160_),
    .ZN(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06719_ (.A1(_01154_),
    .A2(_01161_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06720_ (.A1(_01133_),
    .A2(_01153_),
    .B(_01162_),
    .C(_01055_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06721_ (.A1(_00996_),
    .A2(_01127_),
    .B(_01163_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _06722_ (.A1(_01090_),
    .A2(_00592_),
    .A3(_01092_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06723_ (.I(_01165_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06724_ (.I(_00664_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06725_ (.A1(_00434_),
    .A2(_01167_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06726_ (.I(\as2650.holding_reg[1] ),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06727_ (.A1(_01169_),
    .A2(_00655_),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06728_ (.A1(_05745_),
    .A2(_05782_),
    .B1(_05783_),
    .B2(_05708_),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06729_ (.A1(_01065_),
    .A2(_00989_),
    .B(_01135_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06730_ (.A1(_01171_),
    .A2(_01064_),
    .B(_01172_),
    .C(_01067_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06731_ (.A1(_01169_),
    .A2(_00665_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06732_ (.A1(_01168_),
    .A2(_01170_),
    .B1(_01173_),
    .B2(_01174_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06733_ (.A1(\as2650.holding_reg[1] ),
    .A2(_01168_),
    .A3(_01173_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06734_ (.A1(_00885_),
    .A2(_01176_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06735_ (.I0(_01169_),
    .I1(_00434_),
    .S(_01167_),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06736_ (.A1(_01178_),
    .A2(_01173_),
    .A3(_01174_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06737_ (.I(_01179_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06738_ (.A1(_01173_),
    .A2(_01174_),
    .B(_01178_),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06739_ (.A1(_01180_),
    .A2(_01181_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06740_ (.A1(_00592_),
    .A2(_01175_),
    .A3(_01177_),
    .B1(_01182_),
    .B2(_01082_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06741_ (.A1(_01069_),
    .A2(_01073_),
    .B(_01031_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06742_ (.I(_01072_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06743_ (.A1(_01185_),
    .A2(_01068_),
    .A3(_01070_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06744_ (.A1(_01176_),
    .A2(_01175_),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06745_ (.A1(_01184_),
    .A2(_01186_),
    .B(_01187_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06746_ (.A1(_01184_),
    .A2(_01187_),
    .A3(_01186_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06747_ (.A1(_00885_),
    .A2(_00515_),
    .A3(_01189_),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06748_ (.A1(_01060_),
    .A2(_01073_),
    .B(_01083_),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06749_ (.A1(_01182_),
    .A2(_01191_),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06750_ (.A1(_01188_),
    .A2(_01190_),
    .B1(_01192_),
    .B2(_01058_),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06751_ (.A1(_01166_),
    .A2(_01178_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06752_ (.A1(_01166_),
    .A2(_01183_),
    .A3(_01193_),
    .B(_01194_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06753_ (.I0(_01164_),
    .I1(_01195_),
    .S(_01000_),
    .Z(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06754_ (.I(_01115_),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06755_ (.I0(\as2650.r123[0][1] ),
    .I1(\as2650.r123_2[0][1] ),
    .S(_05710_),
    .Z(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06756_ (.I(_01198_),
    .Z(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06757_ (.I(_01199_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06758_ (.I(_01200_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06759_ (.A1(_01135_),
    .A2(_01021_),
    .A3(_01111_),
    .A4(_01201_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06760_ (.I(_01136_),
    .Z(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06761_ (.I(_01201_),
    .Z(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06762_ (.A1(_01203_),
    .A2(_01112_),
    .B1(_01204_),
    .B2(_01101_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06763_ (.A1(_01202_),
    .A2(_01205_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06764_ (.I(_01106_),
    .Z(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06765_ (.A1(\as2650.r123[1][1] ),
    .A2(_01197_),
    .B1(_01206_),
    .B2(_01207_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06766_ (.A1(_00999_),
    .A2(_01196_),
    .B(_01208_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06767_ (.A1(_01134_),
    .A2(_01200_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06768_ (.I(_05814_),
    .Z(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06769_ (.A1(_01210_),
    .A2(_01111_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06770_ (.I(_01199_),
    .Z(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06771_ (.A1(_05814_),
    .A2(_01134_),
    .A3(_01110_),
    .A4(_01212_),
    .Z(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06772_ (.I(_01213_),
    .Z(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06773_ (.A1(_01209_),
    .A2(_01211_),
    .B(_01214_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06774_ (.I0(\as2650.r123[0][2] ),
    .I1(\as2650.r123_2[0][2] ),
    .S(net51),
    .Z(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06775_ (.I(_01216_),
    .Z(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06776_ (.I(_01217_),
    .Z(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06777_ (.I(_01218_),
    .Z(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06778_ (.A1(_01020_),
    .A2(_01219_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06779_ (.A1(_01215_),
    .A2(_01220_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06780_ (.A1(_01202_),
    .A2(_01221_),
    .Z(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06781_ (.I(_01107_),
    .Z(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06782_ (.A1(\as2650.r123[1][2] ),
    .A2(_01116_),
    .B1(_01222_),
    .B2(_01223_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06783_ (.I(_01114_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06784_ (.I(_00968_),
    .Z(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06785_ (.I(_05757_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06786_ (.I(_01067_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06787_ (.A1(\as2650.holding_reg[2] ),
    .A2(_01228_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06788_ (.A1(_01227_),
    .A2(_01228_),
    .B(_01229_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06789_ (.A1(_01065_),
    .A2(_01064_),
    .B(_01210_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06790_ (.A1(_00421_),
    .A2(_01064_),
    .B(_01231_),
    .C(_00828_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06791_ (.A1(_00423_),
    .A2(_01228_),
    .B(_01232_),
    .C(\as2650.holding_reg[2] ),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06792_ (.I(_01227_),
    .Z(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06793_ (.A1(\as2650.holding_reg[2] ),
    .A2(_00655_),
    .B(_01232_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06794_ (.A1(_01234_),
    .A2(_00829_),
    .B(_01229_),
    .C(_01235_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06795_ (.A1(_01233_),
    .A2(_01236_),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06796_ (.I(_01237_),
    .Z(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06797_ (.A1(_01187_),
    .A2(_01191_),
    .B(_01176_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06798_ (.A1(_01238_),
    .A2(_01239_),
    .B(_00839_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06799_ (.A1(_01238_),
    .A2(_01239_),
    .B(_01240_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06800_ (.A1(_01180_),
    .A2(_01188_),
    .B(_01237_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06801_ (.A1(_01180_),
    .A2(_01188_),
    .A3(_01238_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06802_ (.A1(_01242_),
    .A2(_01243_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06803_ (.I(_01233_),
    .Z(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06804_ (.I(_01245_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06805_ (.A1(_01086_),
    .A2(_01246_),
    .B1(_01236_),
    .B2(_01088_),
    .C(_01165_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06806_ (.A1(_01082_),
    .A2(_01238_),
    .B1(_01244_),
    .B2(_01077_),
    .C(_01247_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06807_ (.A1(_01094_),
    .A2(_01230_),
    .B1(_01241_),
    .B2(_01248_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06808_ (.A1(_00970_),
    .A2(_00987_),
    .A3(_00995_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06809_ (.I(_01250_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _06810_ (.A1(_00430_),
    .A2(_05808_),
    .A3(_05792_),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06811_ (.A1(_01015_),
    .A2(_00432_),
    .B(_01227_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06812_ (.A1(_01252_),
    .A2(_01123_),
    .A3(_01253_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _06813_ (.A1(_00430_),
    .A2(_05808_),
    .A3(_05792_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06814_ (.A1(_01138_),
    .A2(_00432_),
    .B(_01227_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06815_ (.A1(_01008_),
    .A2(_01009_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06816_ (.A1(_01255_),
    .A2(_01256_),
    .B(_01257_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06817_ (.A1(_01257_),
    .A2(_01123_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06818_ (.A1(_00423_),
    .A2(_01259_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06819_ (.A1(_01254_),
    .A2(_01258_),
    .A3(_01260_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06820_ (.I(_01210_),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06821_ (.I(_01262_),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06822_ (.I(_01051_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06823_ (.I(_05766_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06824_ (.A1(_01265_),
    .A2(_01065_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06825_ (.A1(_05745_),
    .A2(_05767_),
    .B1(_05768_),
    .B2(_05739_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06826_ (.A1(_01266_),
    .A2(_01267_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06827_ (.I(_01268_),
    .Z(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06828_ (.A1(_00426_),
    .A2(_01045_),
    .Z(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06829_ (.I(net10),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06830_ (.I(_01271_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06831_ (.I(_01272_),
    .Z(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06832_ (.I(_01273_),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06833_ (.A1(_01274_),
    .A2(_01045_),
    .B(_01036_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06834_ (.A1(_01269_),
    .A2(_01036_),
    .B1(_01270_),
    .B2(_01275_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06835_ (.I(_01034_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06836_ (.A1(_01277_),
    .A2(_01140_),
    .B(_00944_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06837_ (.A1(_01140_),
    .A2(_01276_),
    .B(_01278_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06838_ (.A1(_01263_),
    .A2(_01264_),
    .B(_01014_),
    .C(_01279_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06839_ (.A1(_01252_),
    .A2(_01157_),
    .A3(_01253_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06840_ (.A1(_01016_),
    .A2(_00977_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06841_ (.A1(_01255_),
    .A2(_01256_),
    .B(_01282_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06842_ (.A1(_01282_),
    .A2(_01157_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06843_ (.A1(_01150_),
    .A2(_01284_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06844_ (.A1(_01281_),
    .A2(_01283_),
    .A3(_01285_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06845_ (.A1(_01133_),
    .A2(_01286_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06846_ (.I(_01250_),
    .Z(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06847_ (.A1(_01280_),
    .A2(_01287_),
    .B(_01288_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06848_ (.I(_01103_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06849_ (.I(_00957_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06850_ (.A1(_01290_),
    .A2(_01291_),
    .A3(_00967_),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06851_ (.I(_01292_),
    .Z(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06852_ (.A1(_01251_),
    .A2(_01261_),
    .B(_01289_),
    .C(_01293_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06853_ (.A1(_01226_),
    .A2(_01249_),
    .B(_01294_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06854_ (.A1(_01225_),
    .A2(_01295_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06855_ (.A1(_01224_),
    .A2(_01296_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06856_ (.I(_00437_),
    .Z(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06857_ (.A1(_01268_),
    .A2(_01255_),
    .Z(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06858_ (.I(_01122_),
    .Z(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06859_ (.A1(_00437_),
    .A2(_01252_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06860_ (.A1(_01008_),
    .A2(_01009_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _06861_ (.A1(_01297_),
    .A2(_01010_),
    .B1(_01298_),
    .B2(_01299_),
    .C1(_01300_),
    .C2(_01301_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06862_ (.I(_01302_),
    .Z(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06863_ (.A1(_00709_),
    .A2(_00585_),
    .A3(_00642_),
    .A4(_00906_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06864_ (.A1(_01001_),
    .A2(_00966_),
    .A3(_01128_),
    .A4(_01304_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06865_ (.I(_01265_),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06866_ (.I(_01027_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06867_ (.I(_05807_),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06868_ (.I(_01308_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06869_ (.I(net11),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06870_ (.A1(_00439_),
    .A2(_00932_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06871_ (.A1(_01310_),
    .A2(_00933_),
    .B(_01144_),
    .C(_01311_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06872_ (.A1(_01309_),
    .A2(_01145_),
    .B(_01027_),
    .C(_01312_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06873_ (.A1(_01234_),
    .A2(_01307_),
    .B(_01313_),
    .C(_01051_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06874_ (.A1(_01306_),
    .A2(_01052_),
    .B(_01314_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06875_ (.I(_01156_),
    .Z(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06876_ (.A1(_01316_),
    .A2(_01298_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06877_ (.A1(_01016_),
    .A2(_00977_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06878_ (.I(_01318_),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06879_ (.A1(_01269_),
    .A2(_01284_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06880_ (.A1(_01319_),
    .A2(_01300_),
    .B(_01320_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06881_ (.A1(_01317_),
    .A2(_01321_),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06882_ (.A1(_01305_),
    .A2(_01315_),
    .B1(_01322_),
    .B2(_01154_),
    .C(_01250_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06883_ (.A1(_01251_),
    .A2(_01303_),
    .B(_01323_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06884_ (.A1(\as2650.holding_reg[3] ),
    .A2(_00829_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06885_ (.A1(_00437_),
    .A2(_00656_),
    .B(_01325_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06886_ (.I(_01077_),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06887_ (.I(_05766_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06888_ (.A1(_05727_),
    .A2(_00988_),
    .B(_01328_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06889_ (.A1(_01267_),
    .A2(_00989_),
    .B(_01329_),
    .C(_00654_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06890_ (.A1(\as2650.holding_reg[3] ),
    .A2(_00654_),
    .B(_01330_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06891_ (.A1(_05770_),
    .A2(_00664_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06892_ (.A1(\as2650.holding_reg[3] ),
    .A2(_01167_),
    .B(_01332_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06893_ (.A1(_01331_),
    .A2(_01333_),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06894_ (.I(_01334_),
    .Z(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06895_ (.A1(_01230_),
    .A2(_01235_),
    .B(_01242_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06896_ (.A1(_01335_),
    .A2(_01336_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06897_ (.A1(_01237_),
    .A2(_01239_),
    .B(_01245_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06898_ (.A1(_01335_),
    .A2(_01338_),
    .B(_01058_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06899_ (.A1(_01335_),
    .A2(_01338_),
    .B(_01339_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06900_ (.I(_01086_),
    .Z(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06901_ (.I(_01331_),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06902_ (.A1(_01342_),
    .A2(_01333_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06903_ (.A1(_01342_),
    .A2(_01333_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06904_ (.A1(_00491_),
    .A2(_01091_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06905_ (.A1(_00884_),
    .A2(_01345_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06906_ (.A1(_01081_),
    .A2(_01343_),
    .B(_01346_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06907_ (.A1(_01341_),
    .A2(_01343_),
    .B1(_01344_),
    .B2(_01347_),
    .C(_01165_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06908_ (.A1(_01327_),
    .A2(_01337_),
    .B(_01340_),
    .C(_01348_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06909_ (.A1(_01096_),
    .A2(_01326_),
    .B(_01349_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06910_ (.I0(_01324_),
    .I1(_01350_),
    .S(_01000_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06911_ (.A1(_01202_),
    .A2(_01221_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06912_ (.A1(_01209_),
    .A2(_01211_),
    .B(_01213_),
    .C(_01220_),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06913_ (.A1(_01328_),
    .A2(_01110_),
    .B1(_01212_),
    .B2(_05814_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06914_ (.A1(_01328_),
    .A2(_05752_),
    .A3(_01110_),
    .A4(_01212_),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06915_ (.A1(_01354_),
    .A2(_01355_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06916_ (.I(_05780_),
    .Z(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06917_ (.I0(\as2650.r123[0][3] ),
    .I1(\as2650.r123_2[0][3] ),
    .S(_05709_),
    .Z(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06918_ (.I(_01358_),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06919_ (.I(_01359_),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06920_ (.A1(_01357_),
    .A2(_05775_),
    .A3(_01218_),
    .A4(_01360_),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06921_ (.I(_01359_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06922_ (.I(_01362_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06923_ (.A1(_01134_),
    .A2(_01219_),
    .B1(_01363_),
    .B2(_01020_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06924_ (.A1(_01361_),
    .A2(_01364_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06925_ (.A1(_01356_),
    .A2(_01365_),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06926_ (.A1(_01214_),
    .A2(_01353_),
    .B(_01366_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06927_ (.A1(_01214_),
    .A2(_01353_),
    .A3(_01366_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06928_ (.A1(_01367_),
    .A2(_01368_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06929_ (.A1(_01352_),
    .A2(_01369_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06930_ (.A1(\as2650.r123[1][3] ),
    .A2(_01197_),
    .B1(_01370_),
    .B2(_01207_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06931_ (.A1(_00999_),
    .A2(_01351_),
    .B(_01371_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06932_ (.A1(_01352_),
    .A2(_01369_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06933_ (.A1(_05766_),
    .A2(_01198_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06934_ (.A1(_05760_),
    .A2(_01109_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06935_ (.A1(_01373_),
    .A2(_01361_),
    .A3(_01374_),
    .Z(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06936_ (.A1(_01357_),
    .A2(_01362_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06937_ (.A1(_05752_),
    .A2(_01218_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06938_ (.I0(\as2650.r123[0][4] ),
    .I1(\as2650.r123_2[0][4] ),
    .S(net51),
    .Z(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06939_ (.I(_01378_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06940_ (.I(_01379_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06941_ (.A1(_05776_),
    .A2(_01380_),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06942_ (.A1(_01376_),
    .A2(_01377_),
    .A3(_01381_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06943_ (.A1(_01375_),
    .A2(_01382_),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06944_ (.A1(_01211_),
    .A2(_01373_),
    .B1(_01365_),
    .B2(_01354_),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06945_ (.A1(_01383_),
    .A2(_01384_),
    .Z(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06946_ (.A1(_01367_),
    .A2(_01385_),
    .Z(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06947_ (.A1(_01372_),
    .A2(_01386_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06948_ (.A1(\as2650.r123[1][4] ),
    .A2(_01116_),
    .B1(_01387_),
    .B2(_01223_),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06949_ (.A1(_01237_),
    .A2(_01239_),
    .B1(_01342_),
    .B2(_01333_),
    .C(_01245_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06950_ (.I(_05763_),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06951_ (.A1(_01390_),
    .A2(_01167_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06952_ (.A1(\as2650.holding_reg[4] ),
    .A2(_00665_),
    .B(_01391_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06953_ (.I(_05760_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06954_ (.A1(_01393_),
    .A2(_00962_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06955_ (.A1(_05806_),
    .A2(_00990_),
    .B(_01394_),
    .C(_00828_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06956_ (.A1(\as2650.holding_reg[4] ),
    .A2(_00655_),
    .B(_01395_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06957_ (.A1(_01392_),
    .A2(_01396_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06958_ (.I(_01397_),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06959_ (.A1(_01344_),
    .A2(_01389_),
    .B(_01398_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06960_ (.A1(_01344_),
    .A2(_01398_),
    .A3(_01389_),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06961_ (.A1(_01058_),
    .A2(_01399_),
    .A3(_01400_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06962_ (.A1(_01230_),
    .A2(_01235_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06963_ (.I(_01179_),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06964_ (.A1(_01403_),
    .A2(_01186_),
    .B1(_01230_),
    .B2(_01235_),
    .C(_01181_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06965_ (.A1(_01342_),
    .A2(_01326_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06966_ (.A1(_01402_),
    .A2(_01335_),
    .A3(_01404_),
    .B(_01405_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06967_ (.A1(_01245_),
    .A2(_01236_),
    .B(_01334_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06968_ (.A1(_01180_),
    .A2(_01188_),
    .B(_01407_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06969_ (.A1(_01398_),
    .A2(_01406_),
    .A3(_01408_),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06970_ (.A1(_01406_),
    .A2(_01408_),
    .B(_01397_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06971_ (.A1(_01077_),
    .A2(_01409_),
    .A3(_01410_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06972_ (.I(_01396_),
    .Z(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06973_ (.A1(_01392_),
    .A2(_01412_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06974_ (.A1(_01392_),
    .A2(_01412_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06975_ (.A1(_01086_),
    .A2(_01413_),
    .B1(_01414_),
    .B2(_01088_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06976_ (.I(_01398_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06977_ (.A1(_00885_),
    .A2(_00766_),
    .A3(_01416_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06978_ (.A1(_01094_),
    .A2(_01415_),
    .A3(_01417_),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06979_ (.A1(\as2650.holding_reg[4] ),
    .A2(_00830_),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06980_ (.A1(_01390_),
    .A2(_00764_),
    .B(_01419_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06981_ (.A1(_01401_),
    .A2(_01411_),
    .A3(_01418_),
    .B1(_01420_),
    .B2(_01094_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06982_ (.I(_01421_),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06983_ (.A1(_00430_),
    .A2(_05808_),
    .A3(_00434_),
    .A4(_05770_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06984_ (.A1(_01390_),
    .A2(_01423_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06985_ (.A1(_01308_),
    .A2(_05810_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06986_ (.I(_01301_),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06987_ (.A1(_01309_),
    .A2(_01259_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06988_ (.A1(_01299_),
    .A2(_01424_),
    .B1(_01425_),
    .B2(_01426_),
    .C(_01427_),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06989_ (.I(_01428_),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06990_ (.I(_01393_),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06991_ (.I(_01297_),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06992_ (.I(_05741_),
    .Z(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06993_ (.I(_01432_),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06994_ (.I(net12),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06995_ (.I(_01434_),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06996_ (.I(_01435_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06997_ (.A1(_01436_),
    .A2(_01045_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06998_ (.A1(_05813_),
    .A2(_01147_),
    .B(_01035_),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06999_ (.A1(_01433_),
    .A2(_01036_),
    .B1(_01437_),
    .B2(_01438_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07000_ (.A1(_01307_),
    .A2(_01439_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07001_ (.A1(_01431_),
    .A2(_01307_),
    .B(_01440_),
    .C(_01052_),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07002_ (.A1(_01430_),
    .A2(_01264_),
    .B(_01013_),
    .C(_01441_),
    .ZN(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07003_ (.A1(_01309_),
    .A2(_01284_),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07004_ (.A1(_01316_),
    .A2(_01424_),
    .B1(_01425_),
    .B2(_01318_),
    .C(_01443_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07005_ (.I(_01444_),
    .Z(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07006_ (.A1(_01133_),
    .A2(_01445_),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07007_ (.A1(_01442_),
    .A2(_01446_),
    .B(_01288_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07008_ (.A1(_01251_),
    .A2(_01429_),
    .B(_01447_),
    .C(_01293_),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07009_ (.A1(_01226_),
    .A2(_01422_),
    .B(_01448_),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07010_ (.A1(_01225_),
    .A2(_01449_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07011_ (.A1(_01388_),
    .A2(_01450_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07012_ (.I(_05802_),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07013_ (.A1(_01308_),
    .A2(_01423_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07014_ (.A1(_01451_),
    .A2(_01452_),
    .Z(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07015_ (.A1(_05802_),
    .A2(_05807_),
    .A3(_05810_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07016_ (.A1(_01138_),
    .A2(_05793_),
    .B(_05741_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07017_ (.A1(_01454_),
    .A2(_01455_),
    .ZN(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _07018_ (.A1(_01432_),
    .A2(_01011_),
    .B1(_01453_),
    .B2(_01299_),
    .C1(_01456_),
    .C2(_01426_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07019_ (.I(_01457_),
    .Z(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07020_ (.I(_05733_),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07021_ (.I(_01390_),
    .Z(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07022_ (.A1(_05744_),
    .A2(_05748_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07023_ (.I(_01461_),
    .Z(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07024_ (.A1(_01433_),
    .A2(_05803_),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07025_ (.I(net1),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07026_ (.I(_01464_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07027_ (.I(_01465_),
    .Z(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07028_ (.A1(_01466_),
    .A2(_00933_),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07029_ (.A1(_01463_),
    .A2(_00933_),
    .B(_01035_),
    .C(_01467_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07030_ (.A1(_01462_),
    .A2(_01046_),
    .B(_01039_),
    .C(_01468_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07031_ (.A1(_01460_),
    .A2(_01140_),
    .B(_01469_),
    .C(_00944_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07032_ (.A1(_01459_),
    .A2(_01137_),
    .B(_01470_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07033_ (.A1(_01451_),
    .A2(_01284_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07034_ (.A1(_01316_),
    .A2(_01453_),
    .B1(_01456_),
    .B2(_01319_),
    .C(_01472_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07035_ (.I(_01473_),
    .Z(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07036_ (.A1(_01154_),
    .A2(_01474_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07037_ (.A1(_01154_),
    .A2(_01471_),
    .B(_01475_),
    .C(_00996_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07038_ (.A1(_00996_),
    .A2(_01458_),
    .B(_01476_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07039_ (.I(\as2650.holding_reg[5] ),
    .Z(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07040_ (.A1(_01478_),
    .A2(_00830_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07041_ (.A1(_01432_),
    .A2(_00830_),
    .B(_01479_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07042_ (.A1(_01432_),
    .A2(_00871_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07043_ (.A1(_05733_),
    .A2(_00962_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07044_ (.A1(_05740_),
    .A2(_00991_),
    .B(_01482_),
    .C(_00656_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07045_ (.A1(_01478_),
    .A2(_01481_),
    .A3(_01483_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07046_ (.A1(_01478_),
    .A2(_00667_),
    .B(_01481_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07047_ (.I(_01228_),
    .Z(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07048_ (.A1(\as2650.holding_reg[5] ),
    .A2(_01486_),
    .B(_01483_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07049_ (.I(_01487_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07050_ (.A1(_01485_),
    .A2(_01488_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07051_ (.A1(_01484_),
    .A2(_01489_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07052_ (.A1(_01420_),
    .A2(_01412_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07053_ (.A1(_00500_),
    .A2(_01491_),
    .A3(_01410_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07054_ (.A1(_01490_),
    .A2(_01492_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07055_ (.A1(_01092_),
    .A2(_01493_),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07056_ (.A1(_01413_),
    .A2(_01400_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07057_ (.A1(_01490_),
    .A2(_01495_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07058_ (.A1(_01485_),
    .A2(_01488_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07059_ (.I(_01088_),
    .Z(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07060_ (.A1(_01341_),
    .A2(_01497_),
    .B1(_01489_),
    .B2(_01498_),
    .C(_01166_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07061_ (.A1(_01059_),
    .A2(_01496_),
    .B(_01499_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _07062_ (.A1(_01096_),
    .A2(_01480_),
    .B1(_01494_),
    .B2(_01500_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07063_ (.I0(_01477_),
    .I1(_01501_),
    .S(_00968_),
    .Z(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07064_ (.A1(_01214_),
    .A2(_01353_),
    .B(_01366_),
    .C(_01385_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07065_ (.A1(_01352_),
    .A2(_01369_),
    .A3(_01386_),
    .B(_01503_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07066_ (.A1(_01383_),
    .A2(_01384_),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07067_ (.A1(_01375_),
    .A2(_01382_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07068_ (.A1(_01328_),
    .A2(_01200_),
    .B(_01361_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07069_ (.A1(_01265_),
    .A2(_01200_),
    .A3(_01361_),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07070_ (.A1(_01507_),
    .A2(_01374_),
    .B(_01508_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07071_ (.I(_01379_),
    .Z(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07072_ (.A1(_01357_),
    .A2(_01510_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07073_ (.A1(_05764_),
    .A2(_01217_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07074_ (.A1(_05751_),
    .A2(_01360_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07075_ (.A1(_01511_),
    .A2(_01512_),
    .A3(_01513_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07076_ (.I0(\as2650.r123[0][5] ),
    .I1(\as2650.r123_2[0][5] ),
    .S(_05710_),
    .Z(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07077_ (.I(_01515_),
    .Z(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07078_ (.I(_01516_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07079_ (.I(_01517_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07080_ (.A1(_01020_),
    .A2(_01518_),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07081_ (.A1(_01514_),
    .A2(_01519_),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07082_ (.A1(_05775_),
    .A2(_01362_),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07083_ (.A1(_05781_),
    .A2(_01362_),
    .B1(_01380_),
    .B2(_05775_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _07084_ (.A1(_01521_),
    .A2(_01511_),
    .B1(_01522_),
    .B2(_01377_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07085_ (.A1(_05759_),
    .A2(_01199_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07086_ (.A1(_05732_),
    .A2(_01109_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07087_ (.A1(_01523_),
    .A2(_01524_),
    .A3(_01525_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07088_ (.A1(_01520_),
    .A2(_01526_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07089_ (.A1(_01506_),
    .A2(_01509_),
    .A3(_01527_),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07090_ (.A1(_01505_),
    .A2(_01528_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07091_ (.A1(_01504_),
    .A2(_01529_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07092_ (.A1(\as2650.r123[1][5] ),
    .A2(_01197_),
    .B1(_01530_),
    .B2(_01107_),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07093_ (.A1(_00999_),
    .A2(_01502_),
    .B(_01531_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07094_ (.A1(_01505_),
    .A2(_01528_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07095_ (.A1(_01504_),
    .A2(_01529_),
    .B(_01532_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07096_ (.A1(_01506_),
    .A2(_01527_),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07097_ (.A1(_01506_),
    .A2(_01527_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07098_ (.A1(_01509_),
    .A2(_01534_),
    .B(_01535_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07099_ (.A1(_01393_),
    .A2(_01201_),
    .B(_01523_),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07100_ (.A1(_01393_),
    .A2(_01201_),
    .A3(_01523_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07101_ (.A1(_01537_),
    .A2(_01525_),
    .B(_01538_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07102_ (.A1(_01520_),
    .A2(_01526_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07103_ (.A1(_05776_),
    .A2(_01514_),
    .A3(_01517_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07104_ (.I0(\as2650.r123[0][6] ),
    .I1(\as2650.r123_2[0][6] ),
    .S(_05709_),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07105_ (.I(_01542_),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07106_ (.A1(_05774_),
    .A2(_01543_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07107_ (.A1(_05781_),
    .A2(_01516_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07108_ (.A1(_05780_),
    .A2(_05774_),
    .A3(_01516_),
    .A4(_01543_),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07109_ (.A1(_01544_),
    .A2(_01545_),
    .B(_01546_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07110_ (.A1(_05750_),
    .A2(_01379_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07111_ (.A1(_05758_),
    .A2(_01217_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07112_ (.A1(_05765_),
    .A2(_01359_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07113_ (.A1(_01548_),
    .A2(_01549_),
    .A3(_01550_),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07114_ (.A1(_01547_),
    .A2(_01551_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07115_ (.A1(_05742_),
    .A2(_01108_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07116_ (.A1(_05751_),
    .A2(_01360_),
    .B1(_01510_),
    .B2(_01357_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _07117_ (.A1(_01376_),
    .A2(_01548_),
    .B1(_01554_),
    .B2(_01512_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07118_ (.A1(_05732_),
    .A2(_01199_),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07119_ (.I(_01556_),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07120_ (.A1(_01553_),
    .A2(_01555_),
    .A3(_01557_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07121_ (.A1(_01541_),
    .A2(_01552_),
    .A3(_01558_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07122_ (.A1(_01540_),
    .A2(_01559_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07123_ (.A1(_01539_),
    .A2(_01560_),
    .ZN(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07124_ (.A1(_01533_),
    .A2(_01536_),
    .A3(_01561_),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07125_ (.I(_01562_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07126_ (.A1(\as2650.r123[1][6] ),
    .A2(_01116_),
    .B1(_01563_),
    .B2(_01207_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07127_ (.I(_05797_),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07128_ (.A1(\as2650.holding_reg[6] ),
    .A2(_00829_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07129_ (.A1(_01565_),
    .A2(_01486_),
    .B(_01566_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07130_ (.I(\as2650.holding_reg[6] ),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07131_ (.I(_05743_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07132_ (.A1(_05748_),
    .A2(_00990_),
    .ZN(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07133_ (.A1(_01569_),
    .A2(_00962_),
    .B(_01570_),
    .C(_00666_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07134_ (.A1(_01568_),
    .A2(_00666_),
    .B(_01571_),
    .ZN(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07135_ (.A1(_01572_),
    .A2(_01567_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07136_ (.A1(_01572_),
    .A2(_01567_),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07137_ (.A1(_01573_),
    .A2(_01574_),
    .Z(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07138_ (.I(_01575_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07139_ (.A1(_01413_),
    .A2(_01400_),
    .A3(_01497_),
    .B(_01489_),
    .ZN(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07140_ (.A1(_01576_),
    .A2(_01577_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07141_ (.A1(_01059_),
    .A2(_01578_),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07142_ (.I(_01575_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07143_ (.A1(_01480_),
    .A2(_01487_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07144_ (.A1(_01480_),
    .A2(_01488_),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07145_ (.A1(_01491_),
    .A2(_01410_),
    .A3(_01581_),
    .B(_01582_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07146_ (.A1(_01580_),
    .A2(_01583_),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07147_ (.I(_01574_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07148_ (.A1(_01082_),
    .A2(_01585_),
    .B(_01346_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07149_ (.A1(_01341_),
    .A2(_01585_),
    .B1(_01586_),
    .B2(_01573_),
    .ZN(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07150_ (.A1(_01327_),
    .A2(_01584_),
    .B(_01587_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07151_ (.A1(_01166_),
    .A2(_01567_),
    .B(_01579_),
    .C(_01588_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07152_ (.A1(_05802_),
    .A2(_05807_),
    .A3(_01423_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07153_ (.A1(_01461_),
    .A2(_01590_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07154_ (.A1(_01316_),
    .A2(_01591_),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07155_ (.A1(_05797_),
    .A2(_01454_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07156_ (.A1(_01319_),
    .A2(_01593_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07157_ (.A1(_01565_),
    .A2(_01017_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07158_ (.A1(_01592_),
    .A2(_01594_),
    .A3(_01595_),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07159_ (.I(_01569_),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07160_ (.I(_01597_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07161_ (.I(_01451_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07162_ (.A1(_05716_),
    .A2(_05722_),
    .A3(_05729_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07163_ (.I(_01600_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07164_ (.I(_01601_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07165_ (.A1(_00928_),
    .A2(_00558_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07166_ (.A1(_00488_),
    .A2(_00922_),
    .A3(_01603_),
    .A4(_00974_),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07167_ (.A1(_00942_),
    .A2(_01604_),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07168_ (.A1(_05801_),
    .A2(_01605_),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07169_ (.I(net2),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07170_ (.I(_01607_),
    .Z(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07171_ (.I(_01608_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07172_ (.I(_01609_),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07173_ (.I(_01610_),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07174_ (.A1(_01611_),
    .A2(_01147_),
    .B(_01144_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07175_ (.A1(_01602_),
    .A2(_01145_),
    .B1(_01606_),
    .B2(_01612_),
    .C(_01027_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07176_ (.A1(_01599_),
    .A2(_01307_),
    .B(_01613_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07177_ (.A1(_01264_),
    .A2(_01614_),
    .ZN(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07178_ (.A1(_01598_),
    .A2(_01264_),
    .B(_01014_),
    .C(_01615_),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07179_ (.A1(_01014_),
    .A2(_01596_),
    .B(_01616_),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _07180_ (.A1(_01565_),
    .A2(_01011_),
    .B1(_01591_),
    .B2(_01299_),
    .C1(_01593_),
    .C2(_01426_),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07181_ (.I(_01618_),
    .Z(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07182_ (.A1(_01288_),
    .A2(_01619_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07183_ (.A1(_01055_),
    .A2(_01617_),
    .B(_01620_),
    .C(_01293_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07184_ (.A1(_01226_),
    .A2(_01589_),
    .B(_01621_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07185_ (.A1(_01225_),
    .A2(_01622_),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07186_ (.A1(_01564_),
    .A2(_01623_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07187_ (.A1(_01536_),
    .A2(_01561_),
    .Z(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07188_ (.A1(_01536_),
    .A2(_01561_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07189_ (.A1(_01533_),
    .A2(_01624_),
    .B(_01625_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07190_ (.A1(_01540_),
    .A2(_01559_),
    .Z(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07191_ (.A1(_01539_),
    .A2(_01560_),
    .B(_01627_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07192_ (.A1(_01555_),
    .A2(_01557_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07193_ (.A1(_01555_),
    .A2(_01557_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07194_ (.A1(_01553_),
    .A2(_01629_),
    .B(_01630_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07195_ (.A1(_01541_),
    .A2(_01552_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07196_ (.A1(_01541_),
    .A2(_01552_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07197_ (.A1(_01632_),
    .A2(_01558_),
    .B(_01633_),
    .ZN(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07198_ (.A1(\as2650.r0[3] ),
    .A2(_01378_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07199_ (.A1(_05765_),
    .A2(_01359_),
    .B1(_01510_),
    .B2(_05751_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07200_ (.A1(_01513_),
    .A2(_01635_),
    .B1(_01636_),
    .B2(_01549_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07201_ (.A1(_05742_),
    .A2(_01198_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07202_ (.A1(_01637_),
    .A2(_01638_),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07203_ (.A1(_05723_),
    .A2(_01109_),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07204_ (.A1(_01639_),
    .A2(_01640_),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07205_ (.A1(_01547_),
    .A2(_01551_),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07206_ (.A1(\as2650.r0[5] ),
    .A2(_01216_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07207_ (.A1(\as2650.r0[4] ),
    .A2(_01358_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07208_ (.A1(_01635_),
    .A2(_01643_),
    .A3(_01644_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07209_ (.A1(\as2650.r0[1] ),
    .A2(_01542_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07210_ (.A1(_05750_),
    .A2(_01515_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07211_ (.I0(\as2650.r123[0][7] ),
    .I1(\as2650.r123_2[0][7] ),
    .S(_05709_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07212_ (.I(_01648_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07213_ (.A1(_05774_),
    .A2(_01649_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07214_ (.A1(_01646_),
    .A2(_01647_),
    .A3(_01650_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07215_ (.A1(_01546_),
    .A2(_01645_),
    .A3(_01651_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07216_ (.A1(_01642_),
    .A2(_01652_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07217_ (.A1(_01641_),
    .A2(_01653_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07218_ (.A1(_01634_),
    .A2(_01654_),
    .Z(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07219_ (.A1(_01631_),
    .A2(_01655_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07220_ (.A1(_01628_),
    .A2(_01656_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07221_ (.A1(_01626_),
    .A2(_01657_),
    .Z(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07222_ (.A1(\as2650.r123[1][7] ),
    .A2(_01197_),
    .B1(_01658_),
    .B2(_01207_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07223_ (.A1(_01029_),
    .A2(_00871_),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07224_ (.A1(\as2650.holding_reg[7] ),
    .A2(_01486_),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07225_ (.A1(_01660_),
    .A2(_01661_),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07226_ (.I(_05724_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07227_ (.I(_01663_),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07228_ (.A1(_01664_),
    .A2(_00990_),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07229_ (.A1(_01029_),
    .A2(_00991_),
    .B(_01665_),
    .C(_01486_),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07230_ (.A1(\as2650.holding_reg[7] ),
    .A2(_00871_),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07231_ (.A1(_01666_),
    .A2(_01667_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07232_ (.A1(_01662_),
    .A2(_01668_),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07233_ (.A1(_01662_),
    .A2(_01668_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07234_ (.A1(_01669_),
    .A2(_01670_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07235_ (.A1(_01580_),
    .A2(_01577_),
    .B(_01574_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07236_ (.A1(_01671_),
    .A2(_01672_),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07237_ (.I(_01669_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07238_ (.I(_01670_),
    .Z(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07239_ (.A1(_01674_),
    .A2(_01675_),
    .ZN(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07240_ (.A1(_01568_),
    .A2(_00764_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07241_ (.A1(_01461_),
    .A2(_00764_),
    .B(_01677_),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07242_ (.A1(_01572_),
    .A2(_01678_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07243_ (.A1(_01576_),
    .A2(_01583_),
    .B(_00825_),
    .C(_01679_),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07244_ (.A1(_01676_),
    .A2(_01680_),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07245_ (.I(_01675_),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07246_ (.A1(_01341_),
    .A2(_01674_),
    .B1(_01682_),
    .B2(_01498_),
    .C(_01165_),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _07247_ (.A1(_01059_),
    .A2(_01673_),
    .B1(_01681_),
    .B2(_01092_),
    .C(_01683_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07248_ (.A1(_01096_),
    .A2(_01662_),
    .B(_01684_),
    .ZN(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07249_ (.I(_01685_),
    .Z(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07250_ (.A1(_05797_),
    .A2(_01454_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07251_ (.A1(_01600_),
    .A2(_01687_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07252_ (.A1(_01451_),
    .A2(_01308_),
    .A3(_01461_),
    .A4(_01423_),
    .ZN(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07253_ (.A1(_01600_),
    .A2(_01689_),
    .Z(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07254_ (.A1(_01257_),
    .A2(_01690_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07255_ (.A1(_01601_),
    .A2(_01011_),
    .B1(_01688_),
    .B2(_01426_),
    .C(_01691_),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07256_ (.I(_01692_),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07257_ (.A1(_01282_),
    .A2(_01690_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07258_ (.A1(_01601_),
    .A2(_01017_),
    .B1(_01688_),
    .B2(_01319_),
    .C(_01694_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07259_ (.I(_01695_),
    .Z(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07260_ (.I(_00793_),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07261_ (.A1(_05796_),
    .A2(_01147_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07262_ (.A1(_01697_),
    .A2(_00934_),
    .B(_01145_),
    .C(_01698_),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07263_ (.A1(_01028_),
    .A2(_00427_),
    .B(_01031_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07264_ (.A1(_01046_),
    .A2(_01700_),
    .B(_01040_),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07265_ (.A1(_01462_),
    .A2(_01040_),
    .B1(_01699_),
    .B2(_01701_),
    .C(_00943_),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07266_ (.A1(_01664_),
    .A2(_01137_),
    .B(_01132_),
    .C(_01702_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07267_ (.A1(_01133_),
    .A2(_01696_),
    .B(_01703_),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07268_ (.A1(_01288_),
    .A2(_01704_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07269_ (.A1(_01251_),
    .A2(_01693_),
    .B(_01705_),
    .C(_01293_),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07270_ (.A1(_01226_),
    .A2(_01686_),
    .B(_01706_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07271_ (.A1(_01225_),
    .A2(_01707_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07272_ (.A1(_01659_),
    .A2(_01708_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07273_ (.I(\as2650.r123[0][0] ),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07274_ (.A1(_01290_),
    .A2(_00848_),
    .A3(_01104_),
    .ZN(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07275_ (.A1(_05681_),
    .A2(_05670_),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07276_ (.A1(_00605_),
    .A2(_01711_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07277_ (.A1(_00785_),
    .A2(_00974_),
    .A3(_00963_),
    .A4(_01712_),
    .ZN(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07278_ (.A1(_01103_),
    .A2(_01713_),
    .B(_01052_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07279_ (.A1(_00947_),
    .A2(_00953_),
    .B(_01305_),
    .C(_01007_),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07280_ (.A1(_01605_),
    .A2(_01714_),
    .A3(_01715_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07281_ (.A1(_00838_),
    .A2(_01716_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07282_ (.A1(_05677_),
    .A2(_01710_),
    .A3(_01717_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07283_ (.I(_01718_),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07284_ (.I(_01719_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07285_ (.I(_01099_),
    .ZN(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07286_ (.I(_01717_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07287_ (.A1(_00477_),
    .A2(_00859_),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07288_ (.I(_01723_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07289_ (.I(_01724_),
    .Z(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07290_ (.A1(_01290_),
    .A2(_01725_),
    .A3(_01104_),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07291_ (.I(_01726_),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07292_ (.I(_01727_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07293_ (.I(net48),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07294_ (.A1(net86),
    .A2(_01729_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07295_ (.A1(net70),
    .A2(_01730_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07296_ (.I(_01731_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07297_ (.I(_01732_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07298_ (.I(_01733_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07299_ (.I(_01734_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07300_ (.I(_01730_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07301_ (.I(_01736_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07302_ (.I(_01737_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07303_ (.I(_01738_),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07304_ (.I(_01739_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07305_ (.I(net86),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07306_ (.I(net48),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07307_ (.A1(_01741_),
    .A2(_01742_),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07308_ (.I(_01743_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07309_ (.I(_01744_),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07310_ (.I(_01745_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07311_ (.I(_01746_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07312_ (.A1(\as2650.stack[7][8] ),
    .A2(_01740_),
    .B1(_01747_),
    .B2(\as2650.stack[6][8] ),
    .ZN(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07313_ (.A1(_01741_),
    .A2(_01729_),
    .ZN(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07314_ (.I(_01749_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07315_ (.I(_01750_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07316_ (.I(_01751_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07317_ (.I(_01752_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07318_ (.A1(net86),
    .A2(_01742_),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07319_ (.I(_01754_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07320_ (.I(_01755_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07321_ (.I(_01756_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07322_ (.I(_01757_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07323_ (.A1(\as2650.stack[5][8] ),
    .A2(_01753_),
    .B1(_01758_),
    .B2(\as2650.stack[4][8] ),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07324_ (.A1(_01735_),
    .A2(_01748_),
    .A3(_01759_),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07325_ (.I(_01757_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07326_ (.I(_01752_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07327_ (.A1(\as2650.stack[3][8] ),
    .A2(_01740_),
    .B1(_01761_),
    .B2(\as2650.stack[0][8] ),
    .C1(_01762_),
    .C2(\as2650.stack[1][8] ),
    .ZN(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07328_ (.I(_01732_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07329_ (.I(_01764_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07330_ (.I(_01765_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07331_ (.A1(\as2650.stack[2][8] ),
    .A2(_01747_),
    .B(_01766_),
    .ZN(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07332_ (.I(net70),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07333_ (.A1(_01768_),
    .A2(net73),
    .ZN(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07334_ (.A1(_01736_),
    .A2(_01769_),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07335_ (.I(_01741_),
    .Z(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07336_ (.I(_01742_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07337_ (.A1(_01771_),
    .A2(_01772_),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07338_ (.A1(_01768_),
    .A2(_01773_),
    .B(net73),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07339_ (.A1(_01770_),
    .A2(_01774_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07340_ (.I(_01775_),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07341_ (.I(_01776_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07342_ (.A1(_01763_),
    .A2(_01767_),
    .B(_01777_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07343_ (.I(_01743_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07344_ (.I(_01779_),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07345_ (.I(_01780_),
    .Z(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07346_ (.I(_01781_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07347_ (.A1(\as2650.stack[9][8] ),
    .A2(_01762_),
    .B1(_01761_),
    .B2(\as2650.stack[8][8] ),
    .C1(\as2650.stack[10][8] ),
    .C2(_01782_),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07348_ (.I(_01765_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07349_ (.A1(\as2650.stack[11][8] ),
    .A2(_01740_),
    .B(_01784_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07350_ (.I(_01731_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07351_ (.I(_01786_),
    .Z(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07352_ (.I(_01787_),
    .Z(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07353_ (.I(_01749_),
    .Z(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07354_ (.I(_01789_),
    .Z(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07355_ (.I(_01790_),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07356_ (.A1(\as2650.stack[14][8] ),
    .A2(_01746_),
    .B1(_01791_),
    .B2(\as2650.stack[13][8] ),
    .ZN(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07357_ (.I(_01754_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07358_ (.I(_01793_),
    .Z(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07359_ (.I(_01794_),
    .Z(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07360_ (.A1(\as2650.stack[15][8] ),
    .A2(_01739_),
    .B1(_01795_),
    .B2(\as2650.stack[12][8] ),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07361_ (.A1(_01788_),
    .A2(_01792_),
    .A3(_01796_),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07362_ (.A1(_01783_),
    .A2(_01785_),
    .B(_01797_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07363_ (.I(_01777_),
    .Z(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07364_ (.A1(_01760_),
    .A2(_01778_),
    .B1(_01798_),
    .B2(_01799_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07365_ (.A1(_01105_),
    .A2(_01710_),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07366_ (.I(_01801_),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07367_ (.I(_01726_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07368_ (.A1(_01100_),
    .A2(_01803_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07369_ (.A1(_01728_),
    .A2(_01800_),
    .B(_01802_),
    .C(_01804_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07370_ (.A1(_01721_),
    .A2(_01722_),
    .B(_01719_),
    .C(_01805_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07371_ (.A1(_01709_),
    .A2(_01720_),
    .B(_01806_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07372_ (.I(\as2650.r123[0][1] ),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07373_ (.I(_01196_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07374_ (.I(_01737_),
    .Z(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07375_ (.I(_01809_),
    .Z(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07376_ (.I(_01810_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07377_ (.I(_01781_),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07378_ (.A1(\as2650.stack[7][9] ),
    .A2(_01811_),
    .B1(_01812_),
    .B2(\as2650.stack[6][9] ),
    .ZN(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07379_ (.I(_01750_),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07380_ (.I(_01814_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07381_ (.I(_01815_),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07382_ (.I(_01755_),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07383_ (.I(_01817_),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07384_ (.I(_01818_),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07385_ (.A1(\as2650.stack[5][9] ),
    .A2(_01816_),
    .B1(_01819_),
    .B2(\as2650.stack[4][9] ),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07386_ (.A1(_01766_),
    .A2(_01813_),
    .A3(_01820_),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07387_ (.I(_01779_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07388_ (.I(_01822_),
    .Z(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07389_ (.I(_01823_),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07390_ (.I(_01755_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07391_ (.I(_01825_),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07392_ (.I(_01826_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07393_ (.I(_01750_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07394_ (.I(_01828_),
    .Z(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07395_ (.I(_01829_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07396_ (.A1(\as2650.stack[2][9] ),
    .A2(_01824_),
    .B1(_01827_),
    .B2(\as2650.stack[0][9] ),
    .C1(_01830_),
    .C2(\as2650.stack[1][9] ),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07397_ (.I(_01810_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07398_ (.A1(\as2650.stack[3][9] ),
    .A2(_01832_),
    .B(_01788_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07399_ (.A1(_01831_),
    .A2(_01833_),
    .B(_01777_),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07400_ (.I(_01809_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07401_ (.I(_01835_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07402_ (.A1(\as2650.stack[9][9] ),
    .A2(_01830_),
    .B1(_01827_),
    .B2(\as2650.stack[8][9] ),
    .C1(\as2650.stack[11][9] ),
    .C2(_01836_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07403_ (.A1(\as2650.stack[10][9] ),
    .A2(_01812_),
    .B(_01788_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07404_ (.I(_01738_),
    .Z(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07405_ (.A1(\as2650.stack[15][9] ),
    .A2(_01839_),
    .B1(_01752_),
    .B2(\as2650.stack[13][9] ),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07406_ (.A1(\as2650.stack[14][9] ),
    .A2(_01781_),
    .B1(_01757_),
    .B2(\as2650.stack[12][9] ),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07407_ (.A1(_01765_),
    .A2(_01840_),
    .A3(_01841_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07408_ (.A1(_01837_),
    .A2(_01838_),
    .B(_01842_),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07409_ (.I(_01775_),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07410_ (.I(_01844_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07411_ (.I(_01845_),
    .Z(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07412_ (.A1(_01821_),
    .A2(_01834_),
    .B1(_01843_),
    .B2(_01846_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07413_ (.A1(_01203_),
    .A2(_01803_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07414_ (.I(_01801_),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07415_ (.A1(_01728_),
    .A2(_01847_),
    .B(_01848_),
    .C(_01849_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07416_ (.A1(_01808_),
    .A2(_01722_),
    .B(_01719_),
    .C(_01850_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07417_ (.A1(_01807_),
    .A2(_01720_),
    .B(_01851_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07418_ (.I(\as2650.r123[0][2] ),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07419_ (.I(_01718_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07420_ (.I(_01788_),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07421_ (.I(_01746_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07422_ (.I(_01795_),
    .Z(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07423_ (.A1(\as2650.stack[6][10] ),
    .A2(_01855_),
    .B1(_01856_),
    .B2(\as2650.stack[4][10] ),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07424_ (.I(_01836_),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07425_ (.I(_01791_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07426_ (.A1(\as2650.stack[7][10] ),
    .A2(_01858_),
    .B1(_01859_),
    .B2(\as2650.stack[5][10] ),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07427_ (.A1(_01854_),
    .A2(_01857_),
    .A3(_01860_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07428_ (.I(_01739_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07429_ (.I(_01795_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07430_ (.A1(\as2650.stack[3][10] ),
    .A2(_01862_),
    .B1(_01863_),
    .B2(\as2650.stack[0][10] ),
    .C1(_01753_),
    .C2(\as2650.stack[1][10] ),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07431_ (.I(_01824_),
    .Z(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07432_ (.I(_01734_),
    .Z(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07433_ (.A1(\as2650.stack[2][10] ),
    .A2(_01865_),
    .B(_01866_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07434_ (.A1(_01864_),
    .A2(_01867_),
    .B(_01846_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07435_ (.I(_01791_),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07436_ (.I(_01746_),
    .Z(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07437_ (.A1(\as2650.stack[9][10] ),
    .A2(_01869_),
    .B1(_01758_),
    .B2(\as2650.stack[8][10] ),
    .C1(\as2650.stack[10][10] ),
    .C2(_01870_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07438_ (.I(_01734_),
    .Z(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07439_ (.A1(\as2650.stack[11][10] ),
    .A2(_01858_),
    .B(_01872_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07440_ (.I(_01810_),
    .Z(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07441_ (.I(_01779_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07442_ (.I(_01875_),
    .Z(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07443_ (.I(_01876_),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07444_ (.A1(\as2650.stack[15][10] ),
    .A2(_01874_),
    .B1(_01877_),
    .B2(\as2650.stack[14][10] ),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07445_ (.I(_01818_),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07446_ (.A1(\as2650.stack[13][10] ),
    .A2(_01816_),
    .B1(_01879_),
    .B2(\as2650.stack[12][10] ),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07447_ (.A1(_01784_),
    .A2(_01878_),
    .A3(_01880_),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07448_ (.A1(_01871_),
    .A2(_01873_),
    .B(_01881_),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07449_ (.I(_01777_),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07450_ (.A1(_01861_),
    .A2(_01868_),
    .B1(_01882_),
    .B2(_01883_),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07451_ (.A1(_01263_),
    .A2(_01803_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07452_ (.A1(_01728_),
    .A2(_01884_),
    .B(_01885_),
    .C(_01849_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07453_ (.A1(_01295_),
    .A2(_01722_),
    .B(_01853_),
    .C(_01886_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07454_ (.A1(_01852_),
    .A2(_01720_),
    .B(_01887_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07455_ (.I(\as2650.r123[0][3] ),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07456_ (.I(_01351_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07457_ (.I(_01726_),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07458_ (.A1(\as2650.stack[7][11] ),
    .A2(_01858_),
    .B1(_01859_),
    .B2(\as2650.stack[5][11] ),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07459_ (.A1(\as2650.stack[6][11] ),
    .A2(_01855_),
    .B1(_01856_),
    .B2(\as2650.stack[4][11] ),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07460_ (.A1(_01854_),
    .A2(_01891_),
    .A3(_01892_),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07461_ (.A1(\as2650.stack[3][11] ),
    .A2(_01862_),
    .B1(_01863_),
    .B2(\as2650.stack[0][11] ),
    .C1(_01753_),
    .C2(\as2650.stack[1][11] ),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07462_ (.A1(\as2650.stack[2][11] ),
    .A2(_01865_),
    .B(_01866_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07463_ (.A1(_01894_),
    .A2(_01895_),
    .B(_01846_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07464_ (.A1(\as2650.stack[9][11] ),
    .A2(_01869_),
    .B1(_01758_),
    .B2(\as2650.stack[8][11] ),
    .C1(\as2650.stack[10][11] ),
    .C2(_01747_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07465_ (.A1(\as2650.stack[11][11] ),
    .A2(_01858_),
    .B(_01872_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07466_ (.A1(\as2650.stack[15][11] ),
    .A2(_01874_),
    .B1(_01877_),
    .B2(\as2650.stack[14][11] ),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07467_ (.I(_01815_),
    .Z(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07468_ (.A1(\as2650.stack[13][11] ),
    .A2(_01900_),
    .B1(_01879_),
    .B2(\as2650.stack[12][11] ),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07469_ (.A1(_01784_),
    .A2(_01899_),
    .A3(_01901_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07470_ (.A1(_01897_),
    .A2(_01898_),
    .B(_01902_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07471_ (.A1(_01893_),
    .A2(_01896_),
    .B1(_01903_),
    .B2(_01883_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07472_ (.I(_01306_),
    .Z(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07473_ (.A1(_01905_),
    .A2(_01803_),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07474_ (.A1(_01890_),
    .A2(_01904_),
    .B(_01906_),
    .C(_01849_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07475_ (.A1(_01889_),
    .A2(_01722_),
    .B(_01853_),
    .C(_01907_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07476_ (.A1(_01888_),
    .A2(_01720_),
    .B(_01908_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07477_ (.I(\as2650.r123[0][4] ),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07478_ (.I(_01719_),
    .Z(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07479_ (.I(_01717_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07480_ (.I(_01836_),
    .Z(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07481_ (.A1(\as2650.stack[7][12] ),
    .A2(_01912_),
    .B1(_01855_),
    .B2(\as2650.stack[6][12] ),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07482_ (.I(_01830_),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07483_ (.A1(\as2650.stack[5][12] ),
    .A2(_01914_),
    .B1(_01856_),
    .B2(\as2650.stack[4][12] ),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07484_ (.A1(_01735_),
    .A2(_01913_),
    .A3(_01915_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07485_ (.A1(\as2650.stack[3][12] ),
    .A2(_01862_),
    .B1(_01863_),
    .B2(\as2650.stack[0][12] ),
    .C1(_01753_),
    .C2(\as2650.stack[1][12] ),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07486_ (.A1(\as2650.stack[2][12] ),
    .A2(_01865_),
    .B(_01872_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07487_ (.A1(_01917_),
    .A2(_01918_),
    .B(_01846_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07488_ (.A1(\as2650.stack[9][12] ),
    .A2(_01869_),
    .B1(_01758_),
    .B2(\as2650.stack[8][12] ),
    .C1(\as2650.stack[11][12] ),
    .C2(_01740_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07489_ (.A1(\as2650.stack[10][12] ),
    .A2(_01865_),
    .B(_01872_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07490_ (.A1(\as2650.stack[14][12] ),
    .A2(_01877_),
    .B1(_01879_),
    .B2(\as2650.stack[12][12] ),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07491_ (.A1(\as2650.stack[15][12] ),
    .A2(_01874_),
    .B1(_01900_),
    .B2(\as2650.stack[13][12] ),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07492_ (.A1(_01784_),
    .A2(_01922_),
    .A3(_01923_),
    .Z(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07493_ (.A1(_01920_),
    .A2(_01921_),
    .B(_01924_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07494_ (.A1(_01916_),
    .A2(_01919_),
    .B1(_01925_),
    .B2(_01799_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07495_ (.I(_01430_),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07496_ (.A1(_01927_),
    .A2(_01727_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07497_ (.A1(_01890_),
    .A2(_01926_),
    .B(_01928_),
    .C(_01802_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07498_ (.A1(_01449_),
    .A2(_01911_),
    .B(_01853_),
    .C(_01929_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07499_ (.A1(_01909_),
    .A2(_01910_),
    .B(_01930_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07500_ (.I(\as2650.r123[0][5] ),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07501_ (.I(_01502_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07502_ (.I(_01836_),
    .Z(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07503_ (.I(_01824_),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07504_ (.A1(\as2650.stack[7][13] ),
    .A2(_01933_),
    .B1(_01934_),
    .B2(\as2650.stack[6][13] ),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07505_ (.I(_01830_),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07506_ (.I(_01827_),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07507_ (.A1(\as2650.stack[5][13] ),
    .A2(_01936_),
    .B1(_01937_),
    .B2(\as2650.stack[4][13] ),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07508_ (.A1(_01854_),
    .A2(_01935_),
    .A3(_01938_),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07509_ (.I(_01739_),
    .Z(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07510_ (.I(_01795_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07511_ (.I(_01791_),
    .Z(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07512_ (.A1(\as2650.stack[3][13] ),
    .A2(_01940_),
    .B1(_01941_),
    .B2(\as2650.stack[0][13] ),
    .C1(_01942_),
    .C2(\as2650.stack[1][13] ),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07513_ (.I(_01824_),
    .Z(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07514_ (.A1(\as2650.stack[2][13] ),
    .A2(_01944_),
    .B(_01866_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07515_ (.A1(_01943_),
    .A2(_01945_),
    .B(_01799_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07516_ (.A1(\as2650.stack[9][13] ),
    .A2(_01942_),
    .B1(_01941_),
    .B2(\as2650.stack[8][13] ),
    .C1(\as2650.stack[11][13] ),
    .C2(_01940_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07517_ (.A1(\as2650.stack[10][13] ),
    .A2(_01944_),
    .B(_01866_),
    .ZN(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07518_ (.A1(\as2650.stack[14][13] ),
    .A2(_01812_),
    .B1(_01816_),
    .B2(\as2650.stack[13][13] ),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07519_ (.A1(\as2650.stack[15][13] ),
    .A2(_01832_),
    .B1(_01819_),
    .B2(\as2650.stack[12][13] ),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07520_ (.A1(_01766_),
    .A2(_01949_),
    .A3(_01950_),
    .Z(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07521_ (.A1(_01947_),
    .A2(_01948_),
    .B(_01951_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07522_ (.A1(_01939_),
    .A2(_01946_),
    .B1(_01952_),
    .B2(_01883_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07523_ (.I(_01459_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07524_ (.A1(_01954_),
    .A2(_01727_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07525_ (.A1(_01890_),
    .A2(_01953_),
    .B(_01955_),
    .C(_01802_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07526_ (.A1(_01932_),
    .A2(_01911_),
    .B(_01853_),
    .C(_01956_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07527_ (.A1(_01931_),
    .A2(_01910_),
    .B(_01957_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07528_ (.I(\as2650.r123[0][6] ),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07529_ (.I(_01874_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07530_ (.A1(\as2650.stack[7][14] ),
    .A2(_01959_),
    .B1(_01944_),
    .B2(\as2650.stack[6][14] ),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07531_ (.I(_01900_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07532_ (.I(_01827_),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07533_ (.A1(\as2650.stack[5][14] ),
    .A2(_01961_),
    .B1(_01962_),
    .B2(\as2650.stack[4][14] ),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07534_ (.A1(_01854_),
    .A2(_01960_),
    .A3(_01963_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07535_ (.A1(\as2650.stack[3][14] ),
    .A2(_01912_),
    .B1(_01856_),
    .B2(\as2650.stack[0][14] ),
    .C1(_01859_),
    .C2(\as2650.stack[1][14] ),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07536_ (.A1(\as2650.stack[2][14] ),
    .A2(_01944_),
    .B(_01735_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07537_ (.A1(_01965_),
    .A2(_01966_),
    .B(_01799_),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _07538_ (.A1(\as2650.stack[9][14] ),
    .A2(_01859_),
    .B1(_01941_),
    .B2(\as2650.stack[8][14] ),
    .C1(\as2650.stack[10][14] ),
    .C2(_01870_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07539_ (.A1(\as2650.stack[11][14] ),
    .A2(_01959_),
    .B(_01735_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07540_ (.A1(\as2650.stack[15][14] ),
    .A2(_01832_),
    .B1(_01761_),
    .B2(\as2650.stack[12][14] ),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07541_ (.A1(\as2650.stack[14][14] ),
    .A2(_01782_),
    .B1(_01762_),
    .B2(\as2650.stack[13][14] ),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07542_ (.A1(_01766_),
    .A2(_01970_),
    .A3(_01971_),
    .Z(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07543_ (.A1(_01968_),
    .A2(_01969_),
    .B(_01972_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07544_ (.A1(_01964_),
    .A2(_01967_),
    .B1(_01973_),
    .B2(_01883_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07545_ (.I(_01598_),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07546_ (.A1(_01975_),
    .A2(_01727_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07547_ (.A1(_01890_),
    .A2(_01974_),
    .B(_01976_),
    .C(_01802_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07548_ (.A1(_01622_),
    .A2(_01911_),
    .B(_01718_),
    .C(_01977_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07549_ (.A1(_01958_),
    .A2(_01910_),
    .B(_01978_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07550_ (.I(\as2650.r123[0][7] ),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07551_ (.I(_01664_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07552_ (.A1(_01980_),
    .A2(_01728_),
    .A3(_01849_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07553_ (.A1(_01707_),
    .A2(_01911_),
    .B(_01718_),
    .C(_01981_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07554_ (.A1(_01979_),
    .A2(_01910_),
    .B(_01982_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07555_ (.I(_01030_),
    .Z(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07556_ (.I(_01983_),
    .Z(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07557_ (.I(_01773_),
    .Z(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07558_ (.A1(_00668_),
    .A2(_00855_),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07559_ (.A1(_00605_),
    .A2(_00974_),
    .A3(_01986_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07560_ (.I(_01987_),
    .Z(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07561_ (.I(_01988_),
    .Z(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07562_ (.I(_01768_),
    .Z(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07563_ (.I(_01990_),
    .Z(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07564_ (.I(net73),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07565_ (.I(_01992_),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07566_ (.A1(_01991_),
    .A2(_01993_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07567_ (.I(_01994_),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07568_ (.A1(_01985_),
    .A2(_01989_),
    .A3(_01995_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07569_ (.I(_01996_),
    .Z(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07570_ (.I(_01997_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07571_ (.I(_01991_),
    .Z(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07572_ (.I(_01993_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07573_ (.I(_02000_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07574_ (.I(_01819_),
    .Z(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07575_ (.I(_02002_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07576_ (.I(_00925_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07577_ (.A1(_00554_),
    .A2(_00904_),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07578_ (.A1(_00817_),
    .A2(_02005_),
    .B(_00956_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07579_ (.A1(_00513_),
    .A2(_00626_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07580_ (.I(_01603_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07581_ (.A1(_00518_),
    .A2(_02006_),
    .B1(_02007_),
    .B2(_02008_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07582_ (.A1(_00948_),
    .A2(_00929_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07583_ (.A1(_00878_),
    .A2(_01080_),
    .A3(_05787_),
    .A4(_02010_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07584_ (.I(_00928_),
    .Z(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07585_ (.A1(_00948_),
    .A2(_02012_),
    .A3(_00576_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07586_ (.A1(_01080_),
    .A2(_02013_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07587_ (.A1(_00701_),
    .A2(_02009_),
    .A3(_02011_),
    .B1(_02014_),
    .B2(_00579_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07588_ (.A1(_00568_),
    .A2(\as2650.last_intr ),
    .A3(net75),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07589_ (.A1(_00470_),
    .A2(_02016_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07590_ (.A1(_02004_),
    .A2(_02015_),
    .B(_02017_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07591_ (.I(_01987_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07592_ (.A1(_00861_),
    .A2(_01104_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07593_ (.A1(_02019_),
    .A2(_02020_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07594_ (.A1(_05676_),
    .A2(_02018_),
    .B(_02021_),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07595_ (.I(_02022_),
    .Z(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07596_ (.A1(_01999_),
    .A2(_02001_),
    .A3(_02003_),
    .A4(_02023_),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07597_ (.I(_02024_),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07598_ (.A1(\as2650.stack[13][0] ),
    .A2(_02025_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07599_ (.I(_01771_),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07600_ (.I(_01729_),
    .Z(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07601_ (.A1(_02027_),
    .A2(_02028_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07602_ (.I(_02029_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07603_ (.I(_01994_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07604_ (.A1(_05675_),
    .A2(_02018_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07605_ (.A1(_02019_),
    .A2(_02020_),
    .A3(_02032_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07606_ (.I(_02033_),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07607_ (.A1(_02030_),
    .A2(_02031_),
    .A3(_02034_),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07608_ (.I(_02035_),
    .Z(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07609_ (.I(net90),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07610_ (.I(_02037_),
    .Z(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07611_ (.I(_02038_),
    .ZN(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07612_ (.I(_02021_),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07613_ (.I(_02040_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07614_ (.I(_02040_),
    .Z(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07615_ (.A1(_01100_),
    .A2(_02042_),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07616_ (.A1(_02039_),
    .A2(_02041_),
    .B(_02043_),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07617_ (.I(_02044_),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07618_ (.I(_01996_),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07619_ (.I(_02046_),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07620_ (.A1(_02036_),
    .A2(_02045_),
    .B(_02047_),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07621_ (.A1(_01984_),
    .A2(_01998_),
    .B1(_02026_),
    .B2(_02048_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07622_ (.I(net79),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07623_ (.I(_02049_),
    .Z(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07624_ (.I(_02050_),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07625_ (.I(_02035_),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07626_ (.I(_02052_),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07627_ (.I(net56),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07628_ (.I(_02054_),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07629_ (.I(_02055_),
    .ZN(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07630_ (.I(_02056_),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07631_ (.A1(_01203_),
    .A2(_02042_),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07632_ (.A1(_02057_),
    .A2(_02041_),
    .B(_02058_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07633_ (.I(_02059_),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07634_ (.A1(_02053_),
    .A2(_02060_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07635_ (.I(_02024_),
    .Z(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07636_ (.I(_02046_),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07637_ (.A1(\as2650.stack[13][1] ),
    .A2(_02062_),
    .B(_02063_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07638_ (.A1(_02051_),
    .A2(_01998_),
    .B1(_02061_),
    .B2(_02064_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07639_ (.I(net49),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07640_ (.I(_02065_),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07641_ (.I(_02066_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07642_ (.A1(\as2650.stack[13][2] ),
    .A2(_02025_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07643_ (.I(net89),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07644_ (.I(_02069_),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07645_ (.I(_02070_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07646_ (.A1(_01263_),
    .A2(_02042_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07647_ (.A1(_02071_),
    .A2(_02041_),
    .B(_02072_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07648_ (.I(_02073_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07649_ (.A1(_02036_),
    .A2(_02074_),
    .B(_02063_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07650_ (.A1(_02067_),
    .A2(_01998_),
    .B1(_02068_),
    .B2(_02075_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07651_ (.I(_01028_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07652_ (.I(_02076_),
    .Z(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07653_ (.I(_02077_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07654_ (.A1(\as2650.stack[13][3] ),
    .A2(_02025_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07655_ (.I(net58),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07656_ (.I(_02080_),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07657_ (.I(_02081_),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07658_ (.I(_02040_),
    .Z(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07659_ (.I(_02021_),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07660_ (.A1(_01905_),
    .A2(_02084_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07661_ (.A1(_02082_),
    .A2(_02083_),
    .B(_02085_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07662_ (.I(_02086_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07663_ (.A1(_02036_),
    .A2(_02087_),
    .B(_02063_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07664_ (.A1(_02078_),
    .A2(_01998_),
    .B1(_02079_),
    .B2(_02088_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07665_ (.I(_00940_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07666_ (.I(_02089_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07667_ (.I(_02090_),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07668_ (.I(_02046_),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07669_ (.I(net60),
    .ZN(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07670_ (.I(_02093_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07671_ (.A1(_01927_),
    .A2(_02042_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07672_ (.A1(_02094_),
    .A2(_02041_),
    .B(_02095_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07673_ (.I(_02096_),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07674_ (.A1(_02036_),
    .A2(_02097_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07675_ (.A1(\as2650.stack[13][4] ),
    .A2(_02062_),
    .B(_02063_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07676_ (.A1(_02091_),
    .A2(_02092_),
    .B1(_02098_),
    .B2(_02099_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07677_ (.I(net52),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07678_ (.I(_02100_),
    .Z(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07679_ (.I(_02101_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07680_ (.A1(\as2650.stack[13][5] ),
    .A2(_02025_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07681_ (.I(_02035_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07682_ (.I(net61),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07683_ (.I(_02105_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07684_ (.I(_02106_),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07685_ (.A1(_01954_),
    .A2(_02084_),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07686_ (.A1(_02107_),
    .A2(_02083_),
    .B(_02108_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07687_ (.I(_02109_),
    .Z(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07688_ (.A1(_02104_),
    .A2(_02110_),
    .B(_01997_),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07689_ (.A1(_02102_),
    .A2(_02092_),
    .B1(_02103_),
    .B2(_02111_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07690_ (.I(_05682_),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07691_ (.I(_02112_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07692_ (.A1(\as2650.stack[13][6] ),
    .A2(_02062_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07693_ (.I(net62),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07694_ (.I(_02115_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07695_ (.A1(_01598_),
    .A2(_02084_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07696_ (.A1(_02116_),
    .A2(_02083_),
    .B(_02117_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07697_ (.I(_02118_),
    .Z(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07698_ (.A1(_02104_),
    .A2(_02119_),
    .B(_01997_),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07699_ (.A1(_02113_),
    .A2(_02092_),
    .B1(_02114_),
    .B2(_02120_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07700_ (.I(_05687_),
    .Z(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07701_ (.I(_02121_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07702_ (.A1(\as2650.stack[13][7] ),
    .A2(_02062_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07703_ (.I(_02040_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07704_ (.I(net63),
    .Z(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07705_ (.I(_02125_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07706_ (.A1(_02126_),
    .A2(_02083_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07707_ (.A1(_01980_),
    .A2(_02124_),
    .B(_02127_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07708_ (.I(_02128_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07709_ (.A1(_02104_),
    .A2(_02129_),
    .B(_01997_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07710_ (.A1(_02122_),
    .A2(_02092_),
    .B1(_02123_),
    .B2(_02130_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07711_ (.I(net59),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07712_ (.A1(_02131_),
    .A2(_01772_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07713_ (.I(_02132_),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07714_ (.I(net70),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07715_ (.I(_02134_),
    .Z(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07716_ (.A1(_02135_),
    .A2(_01993_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07717_ (.I(_02136_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07718_ (.I(_01988_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07719_ (.A1(_02133_),
    .A2(_02137_),
    .A3(_02138_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07720_ (.I(_02139_),
    .Z(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07721_ (.I(_02140_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07722_ (.I(_01782_),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07723_ (.I(_02142_),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07724_ (.I(_01993_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07725_ (.A1(_01991_),
    .A2(_02144_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07726_ (.I(_02145_),
    .Z(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07727_ (.I(_02022_),
    .Z(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07728_ (.A1(_02143_),
    .A2(_02146_),
    .A3(_02147_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07729_ (.I(_02148_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07730_ (.A1(\as2650.stack[11][0] ),
    .A2(_02149_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07731_ (.I(_02044_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07732_ (.A1(_02131_),
    .A2(_01729_),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07733_ (.I(_02152_),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07734_ (.I(_02153_),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07735_ (.A1(_02154_),
    .A2(_02137_),
    .A3(_02034_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07736_ (.I(_02155_),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07737_ (.I(_02139_),
    .Z(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07738_ (.I(_02157_),
    .Z(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07739_ (.A1(_02151_),
    .A2(_02156_),
    .B(_02158_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07740_ (.A1(_01984_),
    .A2(_02141_),
    .B1(_02150_),
    .B2(_02159_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07741_ (.I(_02155_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07742_ (.I(_02160_),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07743_ (.A1(_02060_),
    .A2(_02161_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07744_ (.I(_02148_),
    .Z(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07745_ (.I(_02157_),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07746_ (.A1(\as2650.stack[11][1] ),
    .A2(_02163_),
    .B(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07747_ (.A1(_02051_),
    .A2(_02141_),
    .B1(_02162_),
    .B2(_02165_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07748_ (.A1(\as2650.stack[11][2] ),
    .A2(_02149_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07749_ (.I(_02073_),
    .Z(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07750_ (.A1(_02167_),
    .A2(_02156_),
    .B(_02164_),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07751_ (.A1(_02067_),
    .A2(_02141_),
    .B1(_02166_),
    .B2(_02168_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07752_ (.A1(\as2650.stack[11][3] ),
    .A2(_02149_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07753_ (.I(_02086_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07754_ (.A1(_02170_),
    .A2(_02156_),
    .B(_02164_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07755_ (.A1(_02078_),
    .A2(_02141_),
    .B1(_02169_),
    .B2(_02171_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07756_ (.I(_02157_),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07757_ (.A1(\as2650.stack[11][4] ),
    .A2(_02149_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07758_ (.I(_02096_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07759_ (.A1(_02174_),
    .A2(_02156_),
    .B(_02164_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07760_ (.A1(_02091_),
    .A2(_02172_),
    .B1(_02173_),
    .B2(_02175_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07761_ (.A1(\as2650.stack[11][5] ),
    .A2(_02163_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07762_ (.I(_02109_),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07763_ (.I(_02155_),
    .Z(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07764_ (.A1(_02177_),
    .A2(_02178_),
    .B(_02140_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07765_ (.A1(_02102_),
    .A2(_02172_),
    .B1(_02176_),
    .B2(_02179_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07766_ (.A1(\as2650.stack[11][6] ),
    .A2(_02163_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07767_ (.I(_02118_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07768_ (.A1(_02181_),
    .A2(_02178_),
    .B(_02140_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07769_ (.A1(_02113_),
    .A2(_02172_),
    .B1(_02180_),
    .B2(_02182_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07770_ (.A1(\as2650.stack[11][7] ),
    .A2(_02163_),
    .ZN(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07771_ (.I(_02128_),
    .Z(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07772_ (.A1(_02184_),
    .A2(_02178_),
    .B(_02140_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07773_ (.A1(_02122_),
    .A2(_02172_),
    .B1(_02183_),
    .B2(_02185_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07774_ (.I(_02132_),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07775_ (.A1(_02186_),
    .A2(_02031_),
    .A3(_02034_),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07776_ (.I(_02187_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07777_ (.I(_02188_),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07778_ (.I(_02020_),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07779_ (.I(_02190_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07780_ (.I(_02084_),
    .Z(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07781_ (.I(net88),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07782_ (.I(_02193_),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07783_ (.I(_02194_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07784_ (.A1(_01112_),
    .A2(_02191_),
    .B1(_02192_),
    .B2(_02195_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07785_ (.I(_02196_),
    .Z(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07786_ (.I(_02029_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07787_ (.A1(_02198_),
    .A2(_01989_),
    .A3(_01995_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07788_ (.I(_02199_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07789_ (.I(_02200_),
    .Z(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07790_ (.I(_02187_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07791_ (.A1(\as2650.stack[14][8] ),
    .A2(_02202_),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07792_ (.A1(_02189_),
    .A2(_02197_),
    .B(_02201_),
    .C(_02203_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07793_ (.I(net87),
    .Z(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07794_ (.I(_02204_),
    .Z(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07795_ (.A1(_01204_),
    .A2(_02191_),
    .B1(_02192_),
    .B2(_02205_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07796_ (.I(_02206_),
    .Z(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07797_ (.I(_02187_),
    .Z(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07798_ (.A1(\as2650.stack[14][9] ),
    .A2(_02208_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07799_ (.I(_02200_),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07800_ (.A1(_02189_),
    .A2(_02207_),
    .B(_02209_),
    .C(_02210_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07801_ (.I(net66),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07802_ (.I(_02211_),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07803_ (.A1(_01219_),
    .A2(_02191_),
    .B1(_02192_),
    .B2(_02212_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07804_ (.I(_02213_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07805_ (.A1(\as2650.stack[14][10] ),
    .A2(_02208_),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07806_ (.A1(_02189_),
    .A2(_02214_),
    .B(_02215_),
    .C(_02210_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07807_ (.I(net67),
    .Z(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07808_ (.I(_02216_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07809_ (.I(_02217_),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07810_ (.A1(_01363_),
    .A2(_02191_),
    .B1(_02192_),
    .B2(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07811_ (.I(_02219_),
    .Z(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07812_ (.A1(\as2650.stack[14][11] ),
    .A2(_02208_),
    .ZN(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07813_ (.A1(_02189_),
    .A2(_02220_),
    .B(_02221_),
    .C(_02210_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07814_ (.I(_02188_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07815_ (.I(_01380_),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07816_ (.I(net68),
    .Z(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07817_ (.I(_02224_),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07818_ (.A1(_02223_),
    .A2(_02190_),
    .B1(_02124_),
    .B2(_02225_),
    .ZN(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07819_ (.I(_02226_),
    .Z(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07820_ (.A1(\as2650.stack[14][12] ),
    .A2(_02208_),
    .ZN(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07821_ (.A1(_02222_),
    .A2(_02227_),
    .B(_02228_),
    .C(_02210_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07822_ (.I(net69),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07823_ (.A1(_01518_),
    .A2(_02190_),
    .B1(_02124_),
    .B2(_02229_),
    .ZN(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07824_ (.I(_02230_),
    .Z(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07825_ (.A1(\as2650.stack[14][13] ),
    .A2(_02188_),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07826_ (.A1(_02222_),
    .A2(_02231_),
    .B(_02232_),
    .C(_02201_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07827_ (.I(_01543_),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07828_ (.I(_02233_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07829_ (.I(net71),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07830_ (.A1(_02234_),
    .A2(_02190_),
    .B1(_02124_),
    .B2(_02235_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07831_ (.I(_02236_),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07832_ (.A1(\as2650.stack[14][14] ),
    .A2(_02188_),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07833_ (.A1(_02222_),
    .A2(_02237_),
    .B(_02238_),
    .C(_02201_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07834_ (.I(_02052_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07835_ (.A1(\as2650.stack[13][8] ),
    .A2(_02104_),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07836_ (.I(_02046_),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07837_ (.A1(_02239_),
    .A2(_02197_),
    .B(_02240_),
    .C(_02241_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07838_ (.I(_02035_),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07839_ (.A1(\as2650.stack[13][9] ),
    .A2(_02242_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07840_ (.A1(_02239_),
    .A2(_02207_),
    .B(_02243_),
    .C(_02241_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07841_ (.A1(\as2650.stack[13][10] ),
    .A2(_02242_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07842_ (.A1(_02239_),
    .A2(_02214_),
    .B(_02244_),
    .C(_02241_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07843_ (.A1(\as2650.stack[13][11] ),
    .A2(_02242_),
    .ZN(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07844_ (.A1(_02239_),
    .A2(_02220_),
    .B(_02245_),
    .C(_02241_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07845_ (.A1(\as2650.stack[13][12] ),
    .A2(_02242_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07846_ (.A1(_02053_),
    .A2(_02227_),
    .B(_02246_),
    .C(_02047_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07847_ (.A1(\as2650.stack[13][13] ),
    .A2(_02052_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07848_ (.A1(_02053_),
    .A2(_02231_),
    .B(_02247_),
    .C(_02047_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07849_ (.A1(\as2650.stack[13][14] ),
    .A2(_02052_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07850_ (.A1(_02053_),
    .A2(_02237_),
    .B(_02248_),
    .C(_02047_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07851_ (.I(_02033_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07852_ (.A1(_01985_),
    .A2(_02031_),
    .A3(_02249_),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07853_ (.I(_02250_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07854_ (.I(_02251_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07855_ (.A1(\as2650.stack[12][8] ),
    .A2(_02251_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07856_ (.I(_01988_),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07857_ (.A1(_02154_),
    .A2(_02136_),
    .A3(_02254_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07858_ (.I(_02255_),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07859_ (.I(_02256_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07860_ (.A1(_02197_),
    .A2(_02252_),
    .B(_02253_),
    .C(_02257_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07861_ (.I(_02250_),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07862_ (.A1(\as2650.stack[12][9] ),
    .A2(_02258_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07863_ (.A1(_02207_),
    .A2(_02252_),
    .B(_02257_),
    .C(_02259_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07864_ (.I(_02250_),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07865_ (.A1(\as2650.stack[12][10] ),
    .A2(_02260_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07866_ (.A1(_02214_),
    .A2(_02252_),
    .B(_02257_),
    .C(_02261_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07867_ (.A1(\as2650.stack[12][11] ),
    .A2(_02260_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07868_ (.A1(_02220_),
    .A2(_02252_),
    .B(_02257_),
    .C(_02262_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07869_ (.I(_02251_),
    .Z(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07870_ (.I(_02256_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07871_ (.A1(\as2650.stack[12][12] ),
    .A2(_02260_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07872_ (.A1(_02227_),
    .A2(_02263_),
    .B(_02264_),
    .C(_02265_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07873_ (.A1(\as2650.stack[12][13] ),
    .A2(_02260_),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07874_ (.A1(_02231_),
    .A2(_02263_),
    .B(_02264_),
    .C(_02266_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07875_ (.A1(\as2650.stack[12][14] ),
    .A2(_02251_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07876_ (.A1(_02237_),
    .A2(_02263_),
    .B(_02264_),
    .C(_02267_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07877_ (.A1(_02198_),
    .A2(_02136_),
    .A3(_02254_),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07878_ (.I(_02268_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07879_ (.I(_02269_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07880_ (.I(_01762_),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07881_ (.I(_02271_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07882_ (.A1(_02272_),
    .A2(_02146_),
    .A3(_02147_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07883_ (.I(_02273_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07884_ (.A1(\as2650.stack[10][0] ),
    .A2(_02274_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07885_ (.I(_02044_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07886_ (.A1(_02186_),
    .A2(_02137_),
    .A3(_02034_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07887_ (.I(_02277_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07888_ (.I(_02278_),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07889_ (.I(_02268_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07890_ (.I(_02280_),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07891_ (.A1(_02276_),
    .A2(_02279_),
    .B(_02281_),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07892_ (.A1(_01984_),
    .A2(_02270_),
    .B1(_02275_),
    .B2(_02282_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07893_ (.A1(\as2650.stack[10][1] ),
    .A2(_02274_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07894_ (.I(_02059_),
    .Z(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07895_ (.I(_02277_),
    .Z(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07896_ (.I(_02280_),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07897_ (.A1(_02284_),
    .A2(_02285_),
    .B(_02286_),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07898_ (.A1(_02051_),
    .A2(_02270_),
    .B1(_02283_),
    .B2(_02287_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07899_ (.A1(\as2650.stack[10][2] ),
    .A2(_02274_),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07900_ (.A1(_02167_),
    .A2(_02285_),
    .B(_02286_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07901_ (.A1(_02067_),
    .A2(_02270_),
    .B1(_02288_),
    .B2(_02289_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07902_ (.A1(\as2650.stack[10][3] ),
    .A2(_02274_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07903_ (.A1(_02170_),
    .A2(_02285_),
    .B(_02286_),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07904_ (.A1(_02078_),
    .A2(_02270_),
    .B1(_02290_),
    .B2(_02291_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07905_ (.I(_02280_),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07906_ (.I(_02273_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07907_ (.A1(\as2650.stack[10][4] ),
    .A2(_02293_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07908_ (.A1(_02174_),
    .A2(_02285_),
    .B(_02286_),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07909_ (.A1(_02091_),
    .A2(_02292_),
    .B1(_02294_),
    .B2(_02295_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07910_ (.A1(\as2650.stack[10][5] ),
    .A2(_02293_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07911_ (.I(_02277_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07912_ (.A1(_02177_),
    .A2(_02297_),
    .B(_02269_),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07913_ (.A1(_02102_),
    .A2(_02292_),
    .B1(_02296_),
    .B2(_02298_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07914_ (.A1(\as2650.stack[10][6] ),
    .A2(_02293_),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07915_ (.A1(_02181_),
    .A2(_02297_),
    .B(_02269_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07916_ (.A1(_02113_),
    .A2(_02292_),
    .B1(_02299_),
    .B2(_02300_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07917_ (.A1(\as2650.stack[10][7] ),
    .A2(_02293_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07918_ (.I(_02128_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07919_ (.A1(_02302_),
    .A2(_02297_),
    .B(_02269_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07920_ (.A1(_02122_),
    .A2(_02292_),
    .B1(_02301_),
    .B2(_02303_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07921_ (.I(_02160_),
    .Z(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07922_ (.A1(\as2650.stack[11][8] ),
    .A2(_02178_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07923_ (.I(_02157_),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07924_ (.A1(_02304_),
    .A2(_02197_),
    .B(_02305_),
    .C(_02306_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07925_ (.I(_02155_),
    .Z(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07926_ (.A1(\as2650.stack[11][9] ),
    .A2(_02307_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07927_ (.A1(_02304_),
    .A2(_02207_),
    .B(_02308_),
    .C(_02306_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07928_ (.A1(\as2650.stack[11][10] ),
    .A2(_02307_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07929_ (.A1(_02304_),
    .A2(_02214_),
    .B(_02309_),
    .C(_02306_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07930_ (.A1(\as2650.stack[11][11] ),
    .A2(_02307_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07931_ (.A1(_02304_),
    .A2(_02220_),
    .B(_02310_),
    .C(_02306_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07932_ (.A1(\as2650.stack[11][12] ),
    .A2(_02307_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07933_ (.A1(_02161_),
    .A2(_02227_),
    .B(_02311_),
    .C(_02158_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07934_ (.A1(\as2650.stack[11][13] ),
    .A2(_02160_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07935_ (.A1(_02161_),
    .A2(_02231_),
    .B(_02312_),
    .C(_02158_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07936_ (.A1(\as2650.stack[11][14] ),
    .A2(_02160_),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07937_ (.A1(_02161_),
    .A2(_02237_),
    .B(_02313_),
    .C(_02158_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07938_ (.I(_02196_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07939_ (.I(_02278_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07940_ (.A1(\as2650.stack[10][8] ),
    .A2(_02297_),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07941_ (.I(_02280_),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07942_ (.A1(_02314_),
    .A2(_02315_),
    .B(_02316_),
    .C(_02317_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07943_ (.I(_02206_),
    .Z(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07944_ (.I(_02277_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07945_ (.A1(\as2650.stack[10][9] ),
    .A2(_02319_),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07946_ (.A1(_02318_),
    .A2(_02315_),
    .B(_02320_),
    .C(_02317_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07947_ (.I(_02213_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07948_ (.A1(\as2650.stack[10][10] ),
    .A2(_02319_),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07949_ (.A1(_02321_),
    .A2(_02315_),
    .B(_02322_),
    .C(_02317_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07950_ (.I(_02219_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07951_ (.A1(\as2650.stack[10][11] ),
    .A2(_02319_),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07952_ (.A1(_02323_),
    .A2(_02315_),
    .B(_02324_),
    .C(_02317_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07953_ (.I(_02226_),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07954_ (.A1(\as2650.stack[10][12] ),
    .A2(_02319_),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07955_ (.A1(_02325_),
    .A2(_02279_),
    .B(_02326_),
    .C(_02281_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07956_ (.I(_02230_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07957_ (.A1(\as2650.stack[10][13] ),
    .A2(_02278_),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07958_ (.A1(_02327_),
    .A2(_02279_),
    .B(_02328_),
    .C(_02281_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07959_ (.I(_02236_),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07960_ (.A1(\as2650.stack[10][14] ),
    .A2(_02278_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07961_ (.A1(_02329_),
    .A2(_02279_),
    .B(_02330_),
    .C(_02281_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07962_ (.I(_05671_),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07963_ (.I(_02331_),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07964_ (.I(_02008_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07965_ (.I(_02333_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07966_ (.A1(_00503_),
    .A2(_01087_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07967_ (.A1(_00837_),
    .A2(_00464_),
    .A3(_02335_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07968_ (.I(_02336_),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07969_ (.A1(_02334_),
    .A2(_02337_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07970_ (.A1(_02332_),
    .A2(_00853_),
    .B(_02338_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07971_ (.A1(_00938_),
    .A2(_02339_),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07972_ (.I(_00476_),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07973_ (.I(_02341_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07974_ (.A1(_02342_),
    .A2(_00630_),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07975_ (.A1(_00811_),
    .A2(net77),
    .B(_02343_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07976_ (.I(_01663_),
    .Z(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07977_ (.I(_02345_),
    .Z(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07978_ (.I(_02346_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07979_ (.I(_02012_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07980_ (.I(_02348_),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07981_ (.I(_02349_),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07982_ (.I(_02350_),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07983_ (.I(_02351_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07984_ (.A1(_02347_),
    .A2(_02352_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07985_ (.A1(_02338_),
    .A2(_02344_),
    .B1(_02353_),
    .B2(_00853_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07986_ (.A1(net4),
    .A2(_02340_),
    .B1(_02354_),
    .B2(_00938_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07987_ (.A1(_00728_),
    .A2(_02355_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07988_ (.I(_02199_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07989_ (.I(_02356_),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07990_ (.A1(_02151_),
    .A2(_02222_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07991_ (.A1(_01999_),
    .A2(_02000_),
    .A3(_02272_),
    .A4(_02023_),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07992_ (.I(_02359_),
    .Z(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07993_ (.A1(\as2650.stack[14][0] ),
    .A2(_02360_),
    .B(_02201_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07994_ (.A1(_01984_),
    .A2(_02357_),
    .B1(_02358_),
    .B2(_02361_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07995_ (.I(_02359_),
    .Z(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07996_ (.A1(\as2650.stack[14][1] ),
    .A2(_02362_),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07997_ (.I(_02059_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07998_ (.I(_02187_),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07999_ (.I(_02200_),
    .Z(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08000_ (.A1(_02364_),
    .A2(_02365_),
    .B(_02366_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08001_ (.A1(_02051_),
    .A2(_02357_),
    .B1(_02363_),
    .B2(_02367_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08002_ (.I(_02073_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08003_ (.A1(_02368_),
    .A2(_02365_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08004_ (.A1(\as2650.stack[14][2] ),
    .A2(_02360_),
    .B(_02366_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08005_ (.A1(_02067_),
    .A2(_02357_),
    .B1(_02369_),
    .B2(_02370_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08006_ (.A1(\as2650.stack[14][3] ),
    .A2(_02362_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08007_ (.A1(_02170_),
    .A2(_02202_),
    .B(_02366_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08008_ (.A1(_02078_),
    .A2(_02357_),
    .B1(_02371_),
    .B2(_02372_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08009_ (.I(_02200_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08010_ (.A1(\as2650.stack[14][4] ),
    .A2(_02362_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08011_ (.A1(_02174_),
    .A2(_02202_),
    .B(_02366_),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08012_ (.A1(_02091_),
    .A2(_02373_),
    .B1(_02374_),
    .B2(_02375_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08013_ (.I(_02109_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08014_ (.A1(_02376_),
    .A2(_02365_),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08015_ (.A1(\as2650.stack[14][5] ),
    .A2(_02360_),
    .B(_02356_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08016_ (.A1(_02102_),
    .A2(_02373_),
    .B1(_02377_),
    .B2(_02378_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08017_ (.A1(\as2650.stack[14][6] ),
    .A2(_02362_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08018_ (.A1(_02181_),
    .A2(_02202_),
    .B(_02356_),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08019_ (.A1(_02113_),
    .A2(_02373_),
    .B1(_02379_),
    .B2(_02380_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08020_ (.I(_02128_),
    .Z(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08021_ (.A1(_02381_),
    .A2(_02365_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08022_ (.A1(\as2650.stack[14][7] ),
    .A2(_02360_),
    .B(_02356_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08023_ (.A1(_02122_),
    .A2(_02373_),
    .B1(_02382_),
    .B2(_02383_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08024_ (.I(_01983_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08025_ (.I(_02255_),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08026_ (.I(_02385_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08027_ (.I(_01832_),
    .Z(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08028_ (.I(_02387_),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08029_ (.A1(_01999_),
    .A2(_02001_),
    .A3(_02388_),
    .A4(_02023_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08030_ (.I(_02389_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08031_ (.A1(\as2650.stack[12][0] ),
    .A2(_02390_),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08032_ (.I(_02250_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08033_ (.A1(_02276_),
    .A2(_02392_),
    .B(_02264_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08034_ (.A1(_02384_),
    .A2(_02386_),
    .B1(_02391_),
    .B2(_02393_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08035_ (.I(_02050_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08036_ (.A1(_02060_),
    .A2(_02263_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08037_ (.I(_02389_),
    .Z(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08038_ (.I(_02256_),
    .Z(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08039_ (.A1(\as2650.stack[12][1] ),
    .A2(_02396_),
    .B(_02397_),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08040_ (.A1(_02394_),
    .A2(_02386_),
    .B1(_02395_),
    .B2(_02398_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08041_ (.I(_02066_),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08042_ (.A1(\as2650.stack[12][2] ),
    .A2(_02390_),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08043_ (.A1(_02167_),
    .A2(_02392_),
    .B(_02397_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08044_ (.A1(_02399_),
    .A2(_02386_),
    .B1(_02400_),
    .B2(_02401_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08045_ (.I(_02077_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08046_ (.A1(\as2650.stack[12][3] ),
    .A2(_02390_),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08047_ (.A1(_02170_),
    .A2(_02392_),
    .B(_02397_),
    .ZN(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08048_ (.A1(_02402_),
    .A2(_02386_),
    .B1(_02403_),
    .B2(_02404_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08049_ (.I(_02090_),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08050_ (.I(_02256_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08051_ (.A1(\as2650.stack[12][4] ),
    .A2(_02390_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08052_ (.A1(_02174_),
    .A2(_02392_),
    .B(_02397_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08053_ (.A1(_02405_),
    .A2(_02406_),
    .B1(_02407_),
    .B2(_02408_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08054_ (.I(_02101_),
    .Z(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08055_ (.A1(\as2650.stack[12][5] ),
    .A2(_02396_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08056_ (.A1(_02177_),
    .A2(_02258_),
    .B(_02385_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08057_ (.A1(_02409_),
    .A2(_02406_),
    .B1(_02410_),
    .B2(_02411_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08058_ (.I(_02112_),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08059_ (.A1(\as2650.stack[12][6] ),
    .A2(_02396_),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08060_ (.A1(_02181_),
    .A2(_02258_),
    .B(_02385_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08061_ (.A1(_02412_),
    .A2(_02406_),
    .B1(_02413_),
    .B2(_02414_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08062_ (.I(_02121_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08063_ (.A1(\as2650.stack[12][7] ),
    .A2(_02396_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08064_ (.A1(_02302_),
    .A2(_02258_),
    .B(_02385_),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08065_ (.A1(_02415_),
    .A2(_02406_),
    .B1(_02416_),
    .B2(_02417_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08066_ (.A1(_01770_),
    .A2(_02249_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08067_ (.I(_02418_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08068_ (.I(_02419_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08069_ (.A1(\as2650.stack[0][8] ),
    .A2(_02419_),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08070_ (.A1(_02153_),
    .A2(_01989_),
    .A3(_01995_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08071_ (.I(_02422_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08072_ (.I(_02423_),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08073_ (.A1(_02314_),
    .A2(_02420_),
    .B(_02421_),
    .C(_02424_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08074_ (.I(_02418_),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08075_ (.A1(\as2650.stack[0][9] ),
    .A2(_02425_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08076_ (.A1(_02318_),
    .A2(_02420_),
    .B(_02424_),
    .C(_02426_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08077_ (.I(_02418_),
    .Z(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08078_ (.A1(\as2650.stack[0][10] ),
    .A2(_02427_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08079_ (.A1(_02321_),
    .A2(_02420_),
    .B(_02424_),
    .C(_02428_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08080_ (.A1(\as2650.stack[0][11] ),
    .A2(_02427_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08081_ (.A1(_02323_),
    .A2(_02420_),
    .B(_02424_),
    .C(_02429_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08082_ (.I(_02419_),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08083_ (.I(_02423_),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08084_ (.A1(\as2650.stack[0][12] ),
    .A2(_02427_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08085_ (.A1(_02325_),
    .A2(_02430_),
    .B(_02431_),
    .C(_02432_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08086_ (.A1(\as2650.stack[0][13] ),
    .A2(_02427_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08087_ (.A1(_02327_),
    .A2(_02430_),
    .B(_02431_),
    .C(_02433_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08088_ (.A1(\as2650.stack[0][14] ),
    .A2(_02419_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08089_ (.A1(_02329_),
    .A2(_02430_),
    .B(_02431_),
    .C(_02434_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08090_ (.I(_02422_),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08091_ (.I(_02435_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08092_ (.I(_01769_),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08093_ (.I(_02022_),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08094_ (.A1(_02388_),
    .A2(_02437_),
    .A3(_02438_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08095_ (.I(_02439_),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08096_ (.A1(\as2650.stack[0][0] ),
    .A2(_02440_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08097_ (.I(_02418_),
    .Z(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08098_ (.A1(_02276_),
    .A2(_02442_),
    .B(_02431_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08099_ (.A1(_02384_),
    .A2(_02436_),
    .B1(_02441_),
    .B2(_02443_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08100_ (.A1(_02060_),
    .A2(_02430_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08101_ (.I(_02439_),
    .Z(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08102_ (.I(_02423_),
    .Z(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08103_ (.A1(\as2650.stack[0][1] ),
    .A2(_02445_),
    .B(_02446_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08104_ (.A1(_02394_),
    .A2(_02436_),
    .B1(_02444_),
    .B2(_02447_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08105_ (.A1(\as2650.stack[0][2] ),
    .A2(_02440_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08106_ (.I(_02073_),
    .Z(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08107_ (.A1(_02449_),
    .A2(_02442_),
    .B(_02446_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08108_ (.A1(_02399_),
    .A2(_02436_),
    .B1(_02448_),
    .B2(_02450_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08109_ (.A1(\as2650.stack[0][3] ),
    .A2(_02440_),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08110_ (.I(_02086_),
    .Z(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08111_ (.A1(_02452_),
    .A2(_02425_),
    .B(_02446_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08112_ (.A1(_02402_),
    .A2(_02436_),
    .B1(_02451_),
    .B2(_02453_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08113_ (.I(_02423_),
    .Z(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08114_ (.A1(\as2650.stack[0][4] ),
    .A2(_02440_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08115_ (.I(_02096_),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08116_ (.A1(_02456_),
    .A2(_02425_),
    .B(_02446_),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08117_ (.A1(_02405_),
    .A2(_02454_),
    .B1(_02455_),
    .B2(_02457_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08118_ (.A1(_02376_),
    .A2(_02442_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08119_ (.A1(\as2650.stack[0][5] ),
    .A2(_02445_),
    .B(_02435_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08120_ (.A1(_02409_),
    .A2(_02454_),
    .B1(_02458_),
    .B2(_02459_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08121_ (.A1(\as2650.stack[0][6] ),
    .A2(_02445_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08122_ (.I(_02118_),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08123_ (.A1(_02461_),
    .A2(_02425_),
    .B(_02435_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08124_ (.A1(_02412_),
    .A2(_02454_),
    .B1(_02460_),
    .B2(_02462_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08125_ (.A1(_02381_),
    .A2(_02442_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08126_ (.A1(\as2650.stack[0][7] ),
    .A2(_02445_),
    .B(_02435_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08127_ (.A1(_02415_),
    .A2(_02454_),
    .B1(_02463_),
    .B2(_02464_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08128_ (.A1(_01933_),
    .A2(_02145_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08129_ (.A1(_02465_),
    .A2(_02249_),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08130_ (.I(_02466_),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08131_ (.I(_02467_),
    .Z(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08132_ (.A1(\as2650.stack[8][8] ),
    .A2(_02467_),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08133_ (.A1(_01991_),
    .A2(_02144_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08134_ (.I(_02470_),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08135_ (.A1(_02153_),
    .A2(_01989_),
    .A3(_02471_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08136_ (.I(_02472_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08137_ (.I(_02473_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08138_ (.A1(_02314_),
    .A2(_02468_),
    .B(_02469_),
    .C(_02474_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08139_ (.I(_02466_),
    .Z(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08140_ (.A1(\as2650.stack[8][9] ),
    .A2(_02475_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08141_ (.A1(_02318_),
    .A2(_02468_),
    .B(_02474_),
    .C(_02476_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08142_ (.I(_02466_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08143_ (.A1(\as2650.stack[8][10] ),
    .A2(_02477_),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08144_ (.A1(_02321_),
    .A2(_02468_),
    .B(_02474_),
    .C(_02478_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08145_ (.A1(\as2650.stack[8][11] ),
    .A2(_02477_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08146_ (.A1(_02323_),
    .A2(_02468_),
    .B(_02474_),
    .C(_02479_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08147_ (.I(_02467_),
    .Z(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08148_ (.I(_02473_),
    .Z(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08149_ (.A1(\as2650.stack[8][12] ),
    .A2(_02477_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08150_ (.A1(_02325_),
    .A2(_02480_),
    .B(_02481_),
    .C(_02482_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08151_ (.A1(\as2650.stack[8][13] ),
    .A2(_02477_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08152_ (.A1(_02327_),
    .A2(_02480_),
    .B(_02481_),
    .C(_02483_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08153_ (.A1(\as2650.stack[8][14] ),
    .A2(_02467_),
    .ZN(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08154_ (.A1(_02329_),
    .A2(_02480_),
    .B(_02481_),
    .C(_02484_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08155_ (.I(_02033_),
    .Z(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08156_ (.I(_02470_),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08157_ (.A1(_02154_),
    .A2(_02485_),
    .A3(_02486_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08158_ (.I(_02487_),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08159_ (.I(_02488_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08160_ (.A1(\as2650.stack[7][8] ),
    .A2(_02488_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08161_ (.I(_01988_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08162_ (.A1(_02133_),
    .A2(_02491_),
    .A3(_02471_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08163_ (.I(_02492_),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08164_ (.I(_02493_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08165_ (.A1(_02314_),
    .A2(_02489_),
    .B(_02490_),
    .C(_02494_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08166_ (.I(_02487_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08167_ (.A1(\as2650.stack[7][9] ),
    .A2(_02495_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08168_ (.A1(_02318_),
    .A2(_02489_),
    .B(_02494_),
    .C(_02496_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08169_ (.I(_02487_),
    .Z(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08170_ (.A1(\as2650.stack[7][10] ),
    .A2(_02497_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08171_ (.A1(_02321_),
    .A2(_02489_),
    .B(_02494_),
    .C(_02498_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08172_ (.A1(\as2650.stack[7][11] ),
    .A2(_02497_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08173_ (.A1(_02323_),
    .A2(_02489_),
    .B(_02494_),
    .C(_02499_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08174_ (.I(_02488_),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08175_ (.I(_02493_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08176_ (.A1(\as2650.stack[7][12] ),
    .A2(_02497_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08177_ (.A1(_02325_),
    .A2(_02500_),
    .B(_02501_),
    .C(_02502_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08178_ (.A1(\as2650.stack[7][13] ),
    .A2(_02497_),
    .ZN(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08179_ (.A1(_02327_),
    .A2(_02500_),
    .B(_02501_),
    .C(_02503_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08180_ (.A1(\as2650.stack[7][14] ),
    .A2(_02488_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08181_ (.A1(_02329_),
    .A2(_02500_),
    .B(_02501_),
    .C(_02504_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08182_ (.I(_02196_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08183_ (.A1(_02186_),
    .A2(_02485_),
    .A3(_02486_),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08184_ (.I(_02506_),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08185_ (.I(_02507_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08186_ (.A1(\as2650.stack[6][8] ),
    .A2(_02507_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08187_ (.A1(_02198_),
    .A2(_02491_),
    .A3(_02471_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08188_ (.I(_02510_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08189_ (.I(_02511_),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08190_ (.A1(_02505_),
    .A2(_02508_),
    .B(_02509_),
    .C(_02512_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08191_ (.I(_02206_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08192_ (.I(_02506_),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08193_ (.A1(\as2650.stack[6][9] ),
    .A2(_02514_),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08194_ (.A1(_02513_),
    .A2(_02508_),
    .B(_02512_),
    .C(_02515_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08195_ (.I(_02213_),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08196_ (.I(_02506_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08197_ (.A1(\as2650.stack[6][10] ),
    .A2(_02517_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08198_ (.A1(_02516_),
    .A2(_02508_),
    .B(_02512_),
    .C(_02518_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08199_ (.I(_02219_),
    .Z(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08200_ (.A1(\as2650.stack[6][11] ),
    .A2(_02517_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08201_ (.A1(_02519_),
    .A2(_02508_),
    .B(_02512_),
    .C(_02520_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08202_ (.I(_02226_),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08203_ (.I(_02507_),
    .Z(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08204_ (.I(_02511_),
    .Z(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08205_ (.A1(\as2650.stack[6][12] ),
    .A2(_02517_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08206_ (.A1(_02521_),
    .A2(_02522_),
    .B(_02523_),
    .C(_02524_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08207_ (.I(_02230_),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08208_ (.A1(\as2650.stack[6][13] ),
    .A2(_02517_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08209_ (.A1(_02525_),
    .A2(_02522_),
    .B(_02523_),
    .C(_02526_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08210_ (.I(_02236_),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08211_ (.A1(\as2650.stack[6][14] ),
    .A2(_02507_),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08212_ (.A1(_02527_),
    .A2(_02522_),
    .B(_02523_),
    .C(_02528_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08213_ (.A1(_02030_),
    .A2(_02485_),
    .A3(_02486_),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08214_ (.I(_02529_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08215_ (.I(_02530_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08216_ (.A1(\as2650.stack[5][8] ),
    .A2(_02530_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08217_ (.A1(_01985_),
    .A2(_02491_),
    .A3(_02471_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08218_ (.I(_02533_),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08219_ (.I(_02534_),
    .Z(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08220_ (.A1(_02505_),
    .A2(_02531_),
    .B(_02532_),
    .C(_02535_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08221_ (.I(_02529_),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08222_ (.A1(\as2650.stack[5][9] ),
    .A2(_02536_),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08223_ (.A1(_02513_),
    .A2(_02531_),
    .B(_02535_),
    .C(_02537_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08224_ (.I(_02529_),
    .Z(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08225_ (.A1(\as2650.stack[5][10] ),
    .A2(_02538_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08226_ (.A1(_02516_),
    .A2(_02531_),
    .B(_02535_),
    .C(_02539_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08227_ (.A1(\as2650.stack[5][11] ),
    .A2(_02538_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08228_ (.A1(_02519_),
    .A2(_02531_),
    .B(_02535_),
    .C(_02540_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08229_ (.I(_02530_),
    .Z(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08230_ (.I(_02534_),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08231_ (.A1(\as2650.stack[5][12] ),
    .A2(_02538_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08232_ (.A1(_02521_),
    .A2(_02541_),
    .B(_02542_),
    .C(_02543_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08233_ (.A1(\as2650.stack[5][13] ),
    .A2(_02538_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08234_ (.A1(_02525_),
    .A2(_02541_),
    .B(_02542_),
    .C(_02544_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08235_ (.A1(\as2650.stack[5][14] ),
    .A2(_02530_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08236_ (.A1(_02527_),
    .A2(_02541_),
    .B(_02542_),
    .C(_02545_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08237_ (.A1(_00898_),
    .A2(_00615_),
    .ZN(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08238_ (.A1(_00992_),
    .A2(_00734_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08239_ (.A1(_00524_),
    .A2(_00758_),
    .A3(_02547_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08240_ (.A1(_00650_),
    .A2(_02546_),
    .A3(_02548_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08241_ (.A1(_00992_),
    .A2(_00747_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08242_ (.A1(_05698_),
    .A2(_00490_),
    .A3(_00614_),
    .A4(_02550_),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08243_ (.I(\as2650.cycle[8] ),
    .Z(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08244_ (.A1(_02552_),
    .A2(_00483_),
    .B(_00729_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08245_ (.A1(_00743_),
    .A2(_00925_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08246_ (.I(_02554_),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08247_ (.A1(_00459_),
    .A2(_00798_),
    .A3(_00658_),
    .A4(_02555_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08248_ (.A1(_00470_),
    .A2(_00569_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08249_ (.I(_02557_),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08250_ (.A1(_02551_),
    .A2(_02553_),
    .A3(_02556_),
    .A4(_02558_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08251_ (.A1(_00785_),
    .A2(_02549_),
    .B(_02559_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08252_ (.A1(_00605_),
    .A2(_00798_),
    .A3(_00873_),
    .A4(_02555_),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08253_ (.A1(_00472_),
    .A2(_00834_),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08254_ (.A1(_02562_),
    .A2(_00850_),
    .A3(_02550_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08255_ (.A1(_02561_),
    .A2(_02563_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08256_ (.A1(_02560_),
    .A2(_02564_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08257_ (.I(_00506_),
    .Z(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08258_ (.A1(_00557_),
    .A2(_02004_),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08259_ (.I(_02567_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08260_ (.I(_02568_),
    .Z(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08261_ (.I(_00602_),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08262_ (.I(_02570_),
    .Z(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08263_ (.A1(_00645_),
    .A2(_00747_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08264_ (.A1(_00686_),
    .A2(_02572_),
    .ZN(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08265_ (.A1(_05670_),
    .A2(_00735_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08266_ (.A1(_00886_),
    .A2(_00686_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08267_ (.A1(_05698_),
    .A2(_02570_),
    .A3(_02574_),
    .A4(_02575_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08268_ (.A1(_02012_),
    .A2(_00841_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08269_ (.A1(_00734_),
    .A2(_01037_),
    .A3(_02562_),
    .A4(_02577_),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08270_ (.A1(_02571_),
    .A2(_02573_),
    .B(_02576_),
    .C(_02578_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08271_ (.A1(_00483_),
    .A2(_01024_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08272_ (.I(_02580_),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08273_ (.I(_00992_),
    .Z(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08274_ (.A1(_00863_),
    .A2(_02582_),
    .ZN(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08275_ (.A1(_00860_),
    .A2(_02583_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08276_ (.A1(_00659_),
    .A2(_01723_),
    .A3(_02550_),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08277_ (.A1(_02581_),
    .A2(_02584_),
    .B(_02585_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08278_ (.A1(_02566_),
    .A2(_02569_),
    .B(_02579_),
    .C(_02586_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08279_ (.A1(_00660_),
    .A2(_00848_),
    .A3(_02574_),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08280_ (.I(_00873_),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08281_ (.A1(_00850_),
    .A2(_02589_),
    .ZN(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08282_ (.A1(_00852_),
    .A2(_00861_),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08283_ (.I(_00649_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08284_ (.A1(_00506_),
    .A2(_02004_),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08285_ (.A1(_02592_),
    .A2(_02593_),
    .B1(_02567_),
    .B2(_01038_),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08286_ (.A1(_00597_),
    .A2(_00603_),
    .A3(_02573_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08287_ (.A1(_00837_),
    .A2(_00481_),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08288_ (.A1(_05696_),
    .A2(_02335_),
    .A3(_02596_),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08289_ (.A1(_02582_),
    .A2(_02337_),
    .A3(_02597_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08290_ (.I(_02547_),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08291_ (.A1(_00506_),
    .A2(_02599_),
    .A3(_02597_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08292_ (.A1(_00912_),
    .A2(_02595_),
    .A3(_02598_),
    .B1(_02600_),
    .B2(_00753_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _08293_ (.A1(_00735_),
    .A2(_00490_),
    .A3(_00495_),
    .B1(_00501_),
    .B2(_02593_),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08294_ (.A1(_02594_),
    .A2(_02601_),
    .A3(_02602_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08295_ (.A1(_02588_),
    .A2(_02590_),
    .A3(_02591_),
    .B(_02603_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08296_ (.A1(_02565_),
    .A2(_02587_),
    .A3(_02604_),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08297_ (.I(_00749_),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08298_ (.I(_02012_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08299_ (.I(_02607_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08300_ (.A1(_01459_),
    .A2(_02608_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08301_ (.I(net75),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08302_ (.I(_01465_),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08303_ (.I(_02611_),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08304_ (.I(_02612_),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08305_ (.I(_02613_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08306_ (.A1(_02341_),
    .A2(_02336_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08307_ (.I(_02615_),
    .Z(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08308_ (.A1(_02614_),
    .A2(_02616_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08309_ (.I(_02331_),
    .Z(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08310_ (.I(_02618_),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08311_ (.A1(_02610_),
    .A2(_02614_),
    .B(_02617_),
    .C(_02619_),
    .ZN(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08312_ (.I(_02571_),
    .Z(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08313_ (.A1(_02609_),
    .A2(_02620_),
    .B(_02621_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08314_ (.A1(_02606_),
    .A2(_02622_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08315_ (.A1(_02610_),
    .A2(_02605_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08316_ (.I(_00678_),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08317_ (.A1(_02605_),
    .A2(_02623_),
    .B(_02624_),
    .C(_02625_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08318_ (.A1(_01985_),
    .A2(_02485_),
    .A3(_02486_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08319_ (.I(_02626_),
    .Z(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08320_ (.I(_02627_),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08321_ (.A1(\as2650.stack[4][8] ),
    .A2(_02627_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08322_ (.A1(_01934_),
    .A2(_01769_),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08323_ (.A1(_02138_),
    .A2(_02630_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08324_ (.I(_02631_),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08325_ (.I(_02632_),
    .Z(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08326_ (.A1(_02505_),
    .A2(_02628_),
    .B(_02629_),
    .C(_02633_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08327_ (.I(_02626_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08328_ (.A1(\as2650.stack[4][9] ),
    .A2(_02634_),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08329_ (.A1(_02513_),
    .A2(_02628_),
    .B(_02633_),
    .C(_02635_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08330_ (.I(_02626_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08331_ (.A1(\as2650.stack[4][10] ),
    .A2(_02636_),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08332_ (.A1(_02516_),
    .A2(_02628_),
    .B(_02633_),
    .C(_02637_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08333_ (.A1(\as2650.stack[4][11] ),
    .A2(_02636_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08334_ (.A1(_02519_),
    .A2(_02628_),
    .B(_02633_),
    .C(_02638_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08335_ (.I(_02627_),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08336_ (.I(_02632_),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08337_ (.A1(\as2650.stack[4][12] ),
    .A2(_02636_),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08338_ (.A1(_02521_),
    .A2(_02639_),
    .B(_02640_),
    .C(_02641_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08339_ (.A1(\as2650.stack[4][13] ),
    .A2(_02636_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08340_ (.A1(_02525_),
    .A2(_02639_),
    .B(_02640_),
    .C(_02642_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08341_ (.A1(\as2650.stack[4][14] ),
    .A2(_02627_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08342_ (.A1(_02527_),
    .A2(_02639_),
    .B(_02640_),
    .C(_02643_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08343_ (.A1(_02249_),
    .A2(_02630_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08344_ (.I(_02644_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08345_ (.I(_02645_),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08346_ (.A1(\as2650.stack[3][8] ),
    .A2(_02645_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08347_ (.I(_02135_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08348_ (.A1(_02648_),
    .A2(_02144_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08349_ (.A1(_02133_),
    .A2(_02649_),
    .A3(_02254_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08350_ (.I(_02650_),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08351_ (.I(_02651_),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08352_ (.A1(_02505_),
    .A2(_02646_),
    .B(_02647_),
    .C(_02652_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08353_ (.I(_02644_),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08354_ (.A1(\as2650.stack[3][9] ),
    .A2(_02653_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08355_ (.A1(_02513_),
    .A2(_02646_),
    .B(_02652_),
    .C(_02654_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08356_ (.I(_02644_),
    .Z(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08357_ (.A1(\as2650.stack[3][10] ),
    .A2(_02655_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08358_ (.A1(_02516_),
    .A2(_02646_),
    .B(_02652_),
    .C(_02656_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08359_ (.A1(\as2650.stack[3][11] ),
    .A2(_02655_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08360_ (.A1(_02519_),
    .A2(_02646_),
    .B(_02652_),
    .C(_02657_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08361_ (.I(_02645_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08362_ (.I(_02651_),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08363_ (.A1(\as2650.stack[3][12] ),
    .A2(_02655_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08364_ (.A1(_02521_),
    .A2(_02658_),
    .B(_02659_),
    .C(_02660_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08365_ (.A1(\as2650.stack[3][13] ),
    .A2(_02655_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08366_ (.A1(_02525_),
    .A2(_02658_),
    .B(_02659_),
    .C(_02661_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08367_ (.A1(\as2650.stack[3][14] ),
    .A2(_02645_),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08368_ (.A1(_02527_),
    .A2(_02658_),
    .B(_02659_),
    .C(_02662_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08369_ (.I(_02196_),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08370_ (.I(_02033_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08371_ (.A1(_02186_),
    .A2(_02649_),
    .A3(_02664_),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08372_ (.I(_02665_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08373_ (.I(_02666_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08374_ (.A1(\as2650.stack[2][8] ),
    .A2(_02666_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08375_ (.A1(_02198_),
    .A2(_02649_),
    .A3(_02254_),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08376_ (.I(_02669_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08377_ (.I(_02670_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08378_ (.A1(_02663_),
    .A2(_02667_),
    .B(_02668_),
    .C(_02671_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08379_ (.I(_02206_),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08380_ (.I(_02665_),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08381_ (.A1(\as2650.stack[2][9] ),
    .A2(_02673_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08382_ (.A1(_02672_),
    .A2(_02667_),
    .B(_02671_),
    .C(_02674_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08383_ (.I(_02213_),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08384_ (.I(_02665_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08385_ (.A1(\as2650.stack[2][10] ),
    .A2(_02676_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08386_ (.A1(_02675_),
    .A2(_02667_),
    .B(_02671_),
    .C(_02677_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08387_ (.I(_02219_),
    .Z(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08388_ (.A1(\as2650.stack[2][11] ),
    .A2(_02676_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08389_ (.A1(_02678_),
    .A2(_02667_),
    .B(_02671_),
    .C(_02679_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08390_ (.I(_02226_),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08391_ (.I(_02666_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08392_ (.I(_02670_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08393_ (.A1(\as2650.stack[2][12] ),
    .A2(_02676_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08394_ (.A1(_02680_),
    .A2(_02681_),
    .B(_02682_),
    .C(_02683_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08395_ (.I(_02230_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08396_ (.A1(\as2650.stack[2][13] ),
    .A2(_02676_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08397_ (.A1(_02684_),
    .A2(_02681_),
    .B(_02682_),
    .C(_02685_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08398_ (.I(_02236_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08399_ (.A1(\as2650.stack[2][14] ),
    .A2(_02666_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08400_ (.A1(_02686_),
    .A2(_02681_),
    .B(_02682_),
    .C(_02687_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08401_ (.A1(_02030_),
    .A2(_02649_),
    .A3(_02664_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08402_ (.I(_02688_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08403_ (.I(_02689_),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08404_ (.A1(\as2650.stack[1][8] ),
    .A2(_02689_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08405_ (.A1(_01770_),
    .A2(_02138_),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08406_ (.I(_02692_),
    .Z(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08407_ (.I(_02693_),
    .Z(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08408_ (.A1(_02663_),
    .A2(_02690_),
    .B(_02691_),
    .C(_02694_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08409_ (.I(_02688_),
    .Z(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08410_ (.A1(\as2650.stack[1][9] ),
    .A2(_02695_),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08411_ (.A1(_02672_),
    .A2(_02690_),
    .B(_02694_),
    .C(_02696_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08412_ (.I(_02688_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08413_ (.A1(\as2650.stack[1][10] ),
    .A2(_02697_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08414_ (.A1(_02675_),
    .A2(_02690_),
    .B(_02694_),
    .C(_02698_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08415_ (.A1(\as2650.stack[1][11] ),
    .A2(_02697_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08416_ (.A1(_02678_),
    .A2(_02690_),
    .B(_02694_),
    .C(_02699_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08417_ (.I(_02689_),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08418_ (.I(_02693_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08419_ (.A1(\as2650.stack[1][12] ),
    .A2(_02697_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08420_ (.A1(_02680_),
    .A2(_02700_),
    .B(_02701_),
    .C(_02702_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08421_ (.A1(\as2650.stack[1][13] ),
    .A2(_02697_),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08422_ (.A1(_02684_),
    .A2(_02700_),
    .B(_02701_),
    .C(_02703_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08423_ (.A1(\as2650.stack[1][14] ),
    .A2(_02689_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08424_ (.A1(_02686_),
    .A2(_02700_),
    .B(_02701_),
    .C(_02704_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08425_ (.A1(_02154_),
    .A2(_02031_),
    .A3(_02664_),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08426_ (.I(_02705_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08427_ (.I(_02706_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08428_ (.A1(\as2650.stack[15][8] ),
    .A2(_02706_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08429_ (.A1(_02133_),
    .A2(_02491_),
    .A3(_01995_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08430_ (.I(_02709_),
    .Z(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08431_ (.I(_02710_),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08432_ (.A1(_02663_),
    .A2(_02707_),
    .B(_02708_),
    .C(_02711_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08433_ (.I(_02705_),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08434_ (.A1(\as2650.stack[15][9] ),
    .A2(_02712_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08435_ (.A1(_02672_),
    .A2(_02707_),
    .B(_02711_),
    .C(_02713_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08436_ (.I(_02705_),
    .Z(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08437_ (.A1(\as2650.stack[15][10] ),
    .A2(_02714_),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08438_ (.A1(_02675_),
    .A2(_02707_),
    .B(_02711_),
    .C(_02715_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08439_ (.A1(\as2650.stack[15][11] ),
    .A2(_02714_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08440_ (.A1(_02678_),
    .A2(_02707_),
    .B(_02711_),
    .C(_02716_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08441_ (.I(_02706_),
    .Z(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08442_ (.I(_02710_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08443_ (.A1(\as2650.stack[15][12] ),
    .A2(_02714_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08444_ (.A1(_02680_),
    .A2(_02717_),
    .B(_02718_),
    .C(_02719_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08445_ (.A1(\as2650.stack[15][13] ),
    .A2(_02714_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08446_ (.A1(_02684_),
    .A2(_02717_),
    .B(_02718_),
    .C(_02720_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08447_ (.A1(\as2650.stack[15][14] ),
    .A2(_02706_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08448_ (.A1(_02686_),
    .A2(_02717_),
    .B(_02718_),
    .C(_02721_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08449_ (.I(_05670_),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08450_ (.I(_02722_),
    .Z(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08451_ (.I(_01724_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08452_ (.A1(_02723_),
    .A2(_00870_),
    .A3(_02724_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08453_ (.A1(_00879_),
    .A2(_00952_),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08454_ (.I(_00602_),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08455_ (.A1(_02723_),
    .A2(_02726_),
    .A3(_02727_),
    .A4(_00883_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08456_ (.A1(_02725_),
    .A2(_02728_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08457_ (.I(_00948_),
    .Z(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08458_ (.A1(_02730_),
    .A2(_02722_),
    .A3(_01037_),
    .A4(_00834_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08459_ (.I(_02348_),
    .Z(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08460_ (.A1(_02732_),
    .A2(_02727_),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08461_ (.A1(_01026_),
    .A2(_02733_),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08462_ (.A1(_00773_),
    .A2(_00964_),
    .A3(_00982_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08463_ (.A1(_02731_),
    .A2(_02734_),
    .A3(_02735_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08464_ (.I(_00950_),
    .Z(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08465_ (.A1(_02582_),
    .A2(_00542_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08466_ (.A1(_00867_),
    .A2(_02583_),
    .B1(_02738_),
    .B2(_00849_),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08467_ (.I(_00964_),
    .Z(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08468_ (.A1(_05671_),
    .A2(_02740_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08469_ (.A1(_00883_),
    .A2(_00832_),
    .A3(_00855_),
    .A4(_02741_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08470_ (.A1(_00763_),
    .A2(_02742_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08471_ (.A1(_02737_),
    .A2(_02569_),
    .A3(_02739_),
    .A4(_02743_),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08472_ (.I(_05681_),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08473_ (.I(_00952_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08474_ (.I(_00703_),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08475_ (.A1(_02746_),
    .A2(_02747_),
    .A3(_00598_),
    .A4(_00603_),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08476_ (.A1(_02745_),
    .A2(_00886_),
    .A3(_02598_),
    .A4(_02748_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08477_ (.A1(_00898_),
    .A2(_00598_),
    .A3(_00616_),
    .A4(_01130_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08478_ (.A1(_02577_),
    .A2(_02750_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08479_ (.A1(_02566_),
    .A2(_02751_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08480_ (.A1(_00831_),
    .A2(_00768_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08481_ (.A1(_02730_),
    .A2(_02753_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08482_ (.A1(_00952_),
    .A2(_00899_),
    .B1(_01986_),
    .B2(_00606_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08483_ (.A1(_02754_),
    .A2(_02755_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08484_ (.A1(_01143_),
    .A2(_02733_),
    .Z(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08485_ (.A1(_00798_),
    .A2(_00615_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08486_ (.I(_00784_),
    .Z(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08487_ (.A1(_02759_),
    .A2(_01711_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08488_ (.A1(_02758_),
    .A2(_02760_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08489_ (.A1(_00754_),
    .A2(_02761_),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08490_ (.A1(_02756_),
    .A2(_02757_),
    .A3(_02762_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08491_ (.I(_00502_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08492_ (.A1(_02764_),
    .A2(_02726_),
    .A3(_02727_),
    .A4(_02333_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08493_ (.A1(_00833_),
    .A2(_02741_),
    .B(_02765_),
    .C(_02584_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08494_ (.A1(_02752_),
    .A2(_02763_),
    .A3(_02766_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08495_ (.I(_02583_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08496_ (.A1(_02730_),
    .A2(_02341_),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08497_ (.A1(_02348_),
    .A2(_02615_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08498_ (.A1(_02747_),
    .A2(_02337_),
    .A3(_02769_),
    .A4(_02770_),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08499_ (.I(_02008_),
    .Z(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08500_ (.A1(_02341_),
    .A2(_02566_),
    .A3(_02772_),
    .A4(_02337_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08501_ (.A1(_00853_),
    .A2(_02768_),
    .B(_02771_),
    .C(_02773_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08502_ (.A1(_02749_),
    .A2(_02767_),
    .A3(_02774_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08503_ (.A1(_02729_),
    .A2(_02736_),
    .A3(_02744_),
    .A4(_02775_),
    .Z(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08504_ (.I(_00865_),
    .Z(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08505_ (.I(_02777_),
    .Z(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08506_ (.A1(_01770_),
    .A2(_01774_),
    .Z(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08507_ (.I(_02779_),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08508_ (.I(_01736_),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08509_ (.I(_02781_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08510_ (.A1(\as2650.stack[7][6] ),
    .A2(_02782_),
    .B1(_01780_),
    .B2(\as2650.stack[6][6] ),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08511_ (.I(_01749_),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08512_ (.I(_02784_),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08513_ (.A1(\as2650.stack[5][6] ),
    .A2(_02785_),
    .B1(_01756_),
    .B2(\as2650.stack[4][6] ),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08514_ (.A1(_01733_),
    .A2(_02783_),
    .A3(_02786_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08515_ (.A1(_02134_),
    .A2(_01736_),
    .Z(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08516_ (.I(_02788_),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08517_ (.A1(\as2650.stack[3][6] ),
    .A2(_02782_),
    .B1(_01751_),
    .B2(\as2650.stack[1][6] ),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08518_ (.A1(\as2650.stack[2][6] ),
    .A2(_01745_),
    .B1(_01756_),
    .B2(\as2650.stack[0][6] ),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08519_ (.A1(_02789_),
    .A2(_02790_),
    .A3(_02791_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08520_ (.A1(_02780_),
    .A2(_02787_),
    .A3(_02792_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08521_ (.I(_01754_),
    .Z(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08522_ (.I(_02794_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08523_ (.A1(\as2650.stack[9][6] ),
    .A2(_02785_),
    .B1(_02795_),
    .B2(\as2650.stack[8][6] ),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08524_ (.A1(\as2650.stack[11][6] ),
    .A2(_02782_),
    .B1(_01745_),
    .B2(\as2650.stack[10][6] ),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08525_ (.A1(_02789_),
    .A2(_02796_),
    .A3(_02797_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08526_ (.I(_02781_),
    .Z(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08527_ (.A1(\as2650.stack[15][6] ),
    .A2(_02799_),
    .B1(_01745_),
    .B2(\as2650.stack[14][6] ),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08528_ (.A1(\as2650.stack[13][6] ),
    .A2(_02785_),
    .B1(_02795_),
    .B2(\as2650.stack[12][6] ),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08529_ (.A1(_01787_),
    .A2(_02800_),
    .A3(_02801_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08530_ (.A1(_01776_),
    .A2(_02798_),
    .A3(_02802_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08531_ (.A1(_02793_),
    .A2(_02803_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08532_ (.I(_02777_),
    .Z(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08533_ (.I(_00878_),
    .Z(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08534_ (.I(_02806_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08535_ (.I(_02807_),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08536_ (.I(_02808_),
    .Z(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08537_ (.I(_02764_),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08538_ (.I(_02810_),
    .Z(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08539_ (.I(_02592_),
    .Z(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08540_ (.I(_02812_),
    .Z(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08541_ (.I(_01037_),
    .Z(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08542_ (.I(_02814_),
    .Z(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08543_ (.A1(_02815_),
    .A2(_01032_),
    .A3(_01454_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08544_ (.A1(_01462_),
    .A2(_02815_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08545_ (.I(_00613_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08546_ (.I(_02818_),
    .Z(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08547_ (.A1(_01597_),
    .A2(_01459_),
    .A3(_01430_),
    .A4(_01265_),
    .Z(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08548_ (.A1(_01210_),
    .A2(_01135_),
    .A3(_01021_),
    .A4(_02820_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08549_ (.A1(_02345_),
    .A2(_02821_),
    .B(_02590_),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08550_ (.I(_02607_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08551_ (.I(_02823_),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08552_ (.A1(_01598_),
    .A2(_02590_),
    .B(_02822_),
    .C(_02824_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08553_ (.I(_01610_),
    .Z(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08554_ (.I(_02596_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08555_ (.A1(net94),
    .A2(_02826_),
    .B(_02723_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08556_ (.A1(_02342_),
    .A2(_02826_),
    .B(_02827_),
    .C(_02828_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08557_ (.A1(_02807_),
    .A2(_01498_),
    .A3(_02829_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08558_ (.A1(_02819_),
    .A2(_02825_),
    .A3(_02830_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08559_ (.A1(_02813_),
    .A2(_02816_),
    .A3(_02817_),
    .A4(_02831_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08560_ (.I(_00594_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08561_ (.I(_01602_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08562_ (.I(_01433_),
    .Z(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08563_ (.I(_01565_),
    .Z(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08564_ (.I(_02836_),
    .Z(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08565_ (.A1(_02834_),
    .A2(_02835_),
    .A3(_05793_),
    .A4(_02837_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08566_ (.A1(_02833_),
    .A2(_01700_),
    .A3(_02838_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08567_ (.A1(_02811_),
    .A2(_02832_),
    .A3(_02839_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08568_ (.I(_00923_),
    .Z(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08569_ (.I(_02841_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08570_ (.A1(_00630_),
    .A2(_02842_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08571_ (.I(_01043_),
    .Z(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08572_ (.I(_02844_),
    .Z(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08573_ (.I(_01142_),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08574_ (.I(_02846_),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08575_ (.I(_01271_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08576_ (.I(_02848_),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08577_ (.I(_02849_),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08578_ (.I(_02850_),
    .Z(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08579_ (.I(net11),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08580_ (.I(_02852_),
    .Z(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08581_ (.I(_02853_),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08582_ (.I(_02854_),
    .Z(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08583_ (.I(_02855_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08584_ (.A1(_02845_),
    .A2(_02847_),
    .A3(_02851_),
    .A4(_02856_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08585_ (.I(_01436_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08586_ (.I(_02858_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08587_ (.I(_02859_),
    .Z(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08588_ (.I(_02826_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08589_ (.A1(_02860_),
    .A2(_02613_),
    .A3(_02861_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08590_ (.A1(_02842_),
    .A2(_02857_),
    .A3(_02862_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08591_ (.A1(_02809_),
    .A2(_02840_),
    .A3(_02843_),
    .A4(_02863_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08592_ (.I(_02722_),
    .Z(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08593_ (.A1(_00880_),
    .A2(_02865_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08594_ (.I(_02866_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08595_ (.A1(_02834_),
    .A2(_00769_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08596_ (.A1(_02346_),
    .A2(_00769_),
    .A3(_02821_),
    .B1(_02868_),
    .B2(_01687_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08597_ (.A1(_02867_),
    .A2(_02869_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08598_ (.A1(_02805_),
    .A2(_02864_),
    .A3(_02870_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08599_ (.A1(net79),
    .A2(_01671_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08600_ (.A1(_01572_),
    .A2(_01678_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08601_ (.A1(_01660_),
    .A2(_01661_),
    .Z(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08602_ (.A1(_02874_),
    .A2(_01668_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08603_ (.A1(_01576_),
    .A2(_01676_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08604_ (.A1(_01420_),
    .A2(_01412_),
    .B1(_01480_),
    .B2(_01488_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08605_ (.A1(_01406_),
    .A2(_01490_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08606_ (.A1(_01581_),
    .A2(_02877_),
    .B1(_02878_),
    .B2(_01416_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08607_ (.A1(_02874_),
    .A2(_01668_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08608_ (.A1(_02873_),
    .A2(_02875_),
    .B1(_02876_),
    .B2(_02879_),
    .C(_02880_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08609_ (.A1(_02872_),
    .A2(_02881_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08610_ (.A1(_02872_),
    .A2(_02881_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08611_ (.A1(_00886_),
    .A2(_00461_),
    .A3(_02883_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08612_ (.A1(_02882_),
    .A2(_02884_),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08613_ (.A1(_01097_),
    .A2(_01195_),
    .A3(_01249_),
    .A4(_01350_),
    .Z(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08614_ (.A1(_01422_),
    .A2(_01501_),
    .A3(_01589_),
    .A4(_02886_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08615_ (.A1(_00958_),
    .A2(_01686_),
    .A3(_02887_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08616_ (.I(_01711_),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08617_ (.I(_02889_),
    .Z(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08618_ (.A1(_02885_),
    .A2(_02888_),
    .B(_02890_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08619_ (.A1(_02778_),
    .A2(_02804_),
    .B1(_02871_),
    .B2(_02891_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08620_ (.I(_00677_),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08621_ (.I(_02893_),
    .Z(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08622_ (.A1(net94),
    .A2(_02776_),
    .B(_02894_),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08623_ (.A1(_02776_),
    .A2(_02892_),
    .B(_02895_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08624_ (.A1(_02347_),
    .A2(_00769_),
    .B(_02868_),
    .C(_02352_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08625_ (.I(_02896_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08626_ (.A1(_01484_),
    .A2(_01489_),
    .B(_01074_),
    .C(_01416_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08627_ (.A1(_01182_),
    .A2(_01407_),
    .A3(_02876_),
    .A4(_02898_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08628_ (.A1(_02882_),
    .A2(_02899_),
    .B(_02884_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08629_ (.I(_02823_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08630_ (.I(_02901_),
    .Z(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08631_ (.I(_02902_),
    .Z(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08632_ (.A1(_00958_),
    .A2(_01686_),
    .B(_02900_),
    .C(_02903_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08633_ (.A1(_02897_),
    .A2(_02904_),
    .B(_00647_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08634_ (.I(_01732_),
    .Z(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08635_ (.I(_02906_),
    .Z(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08636_ (.I(_02781_),
    .Z(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08637_ (.I(_01822_),
    .Z(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08638_ (.A1(\as2650.stack[7][7] ),
    .A2(_02908_),
    .B1(_02909_),
    .B2(\as2650.stack[6][7] ),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08639_ (.A1(\as2650.stack[5][7] ),
    .A2(_01790_),
    .B1(_01794_),
    .B2(\as2650.stack[4][7] ),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08640_ (.A1(_02907_),
    .A2(_02910_),
    .A3(_02911_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08641_ (.I(_02784_),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08642_ (.I(_02794_),
    .Z(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08643_ (.A1(\as2650.stack[1][7] ),
    .A2(_02913_),
    .B1(_02914_),
    .B2(\as2650.stack[0][7] ),
    .C1(\as2650.stack[3][7] ),
    .C2(_02799_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08644_ (.A1(\as2650.stack[2][7] ),
    .A2(_02909_),
    .B(_01733_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08645_ (.A1(_02915_),
    .A2(_02916_),
    .B(_01844_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08646_ (.A1(\as2650.stack[9][7] ),
    .A2(_02913_),
    .B1(_02795_),
    .B2(\as2650.stack[8][7] ),
    .C1(\as2650.stack[11][7] ),
    .C2(_02799_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08647_ (.A1(\as2650.stack[10][7] ),
    .A2(_02909_),
    .B(_01764_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08648_ (.A1(\as2650.stack[14][7] ),
    .A2(_01875_),
    .B1(_01817_),
    .B2(\as2650.stack[12][7] ),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08649_ (.A1(\as2650.stack[15][7] ),
    .A2(_01809_),
    .B1(_01814_),
    .B2(\as2650.stack[13][7] ),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08650_ (.A1(_01764_),
    .A2(_02920_),
    .A3(_02921_),
    .Z(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08651_ (.A1(_02918_),
    .A2(_02919_),
    .B(_02922_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08652_ (.A1(_02912_),
    .A2(_02917_),
    .B1(_02923_),
    .B2(_01845_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08653_ (.A1(_02805_),
    .A2(_02924_),
    .B(_02776_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08654_ (.A1(_00843_),
    .A2(_01090_),
    .A3(_00493_),
    .A4(_00464_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08655_ (.I(net74),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08656_ (.A1(_02135_),
    .A2(_02849_),
    .B1(_01436_),
    .B2(_02927_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08657_ (.A1(_01772_),
    .A2(_01043_),
    .B1(_01142_),
    .B2(_01771_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08658_ (.I(net85),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08659_ (.I(net77),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08660_ (.I(_00792_),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08661_ (.I(net1),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08662_ (.A1(_01992_),
    .A2(_01310_),
    .B1(_02933_),
    .B2(_02610_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08663_ (.A1(_02930_),
    .A2(_01611_),
    .B1(_02931_),
    .B2(_02932_),
    .C(_02934_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08664_ (.A1(_02928_),
    .A2(_02929_),
    .A3(_02935_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08665_ (.A1(_02342_),
    .A2(_02335_),
    .A3(_02827_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08666_ (.A1(_05695_),
    .A2(_00493_),
    .A3(_02827_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08667_ (.A1(_05687_),
    .A2(_00792_),
    .B1(_01042_),
    .B2(_01030_),
    .C1(_02076_),
    .C2(_02854_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08668_ (.I(_01608_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08669_ (.A1(_02049_),
    .A2(_01141_),
    .B1(_01466_),
    .B2(_02100_),
    .C1(_02940_),
    .C2(_05682_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08670_ (.A1(_02065_),
    .A2(_02848_),
    .B1(_01435_),
    .B2(_02089_),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08671_ (.A1(_02939_),
    .A2(_02941_),
    .A3(_02942_),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08672_ (.A1(_01141_),
    .A2(_01034_),
    .B1(_01297_),
    .B2(_02853_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08673_ (.A1(_02848_),
    .A2(_01234_),
    .B1(_02836_),
    .B2(_02940_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08674_ (.A1(_00626_),
    .A2(_01601_),
    .B1(_01138_),
    .B2(_01042_),
    .C1(_01460_),
    .C2(_01435_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08675_ (.A1(_02944_),
    .A2(_02945_),
    .A3(_02946_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08676_ (.A1(_01466_),
    .A2(_01433_),
    .B(_02938_),
    .C(_02947_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08677_ (.A1(_02938_),
    .A2(_02943_),
    .B(_02926_),
    .C(_02948_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08678_ (.A1(_02926_),
    .A2(_02936_),
    .B(_02937_),
    .C(_02949_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08679_ (.I(net54),
    .Z(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08680_ (.I(_02932_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08681_ (.A1(_02951_),
    .A2(_02952_),
    .A3(_02335_),
    .A4(_02827_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08682_ (.A1(_02597_),
    .A2(_02950_),
    .A3(_02953_),
    .Z(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08683_ (.I(_01697_),
    .Z(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08684_ (.I(_02597_),
    .Z(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08685_ (.A1(_02951_),
    .A2(_02955_),
    .A3(_02956_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08686_ (.A1(_02954_),
    .A2(_02957_),
    .B(_02351_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08687_ (.A1(_02346_),
    .A2(_02902_),
    .B(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08688_ (.I(_02592_),
    .Z(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08689_ (.A1(_02960_),
    .A2(_01700_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08690_ (.A1(_00951_),
    .A2(_02959_),
    .B(_02961_),
    .C(_02817_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08691_ (.A1(_02811_),
    .A2(_02962_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08692_ (.A1(_00865_),
    .A2(_02807_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08693_ (.I(_02964_),
    .Z(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08694_ (.A1(_02843_),
    .A2(_02963_),
    .B(_02965_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08695_ (.A1(_02925_),
    .A2(_02966_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08696_ (.A1(_02951_),
    .A2(_02776_),
    .B(_02894_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08697_ (.A1(_02905_),
    .A2(_02967_),
    .B(_02968_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08698_ (.I(_02709_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08699_ (.I(_02969_),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08700_ (.A1(_01999_),
    .A2(_02001_),
    .A3(_02143_),
    .A4(_02023_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08701_ (.I(_02971_),
    .Z(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08702_ (.A1(\as2650.stack[15][0] ),
    .A2(_02972_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08703_ (.I(_02705_),
    .Z(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08704_ (.A1(_02276_),
    .A2(_02974_),
    .B(_02718_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08705_ (.A1(_02384_),
    .A2(_02970_),
    .B1(_02973_),
    .B2(_02975_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08706_ (.I(_02059_),
    .Z(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08707_ (.A1(_02976_),
    .A2(_02717_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08708_ (.I(_02971_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08709_ (.I(_02710_),
    .Z(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08710_ (.A1(\as2650.stack[15][1] ),
    .A2(_02978_),
    .B(_02979_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08711_ (.A1(_02394_),
    .A2(_02970_),
    .B1(_02977_),
    .B2(_02980_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08712_ (.A1(\as2650.stack[15][2] ),
    .A2(_02972_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08713_ (.A1(_02449_),
    .A2(_02974_),
    .B(_02979_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08714_ (.A1(_02399_),
    .A2(_02970_),
    .B1(_02981_),
    .B2(_02982_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08715_ (.A1(\as2650.stack[15][3] ),
    .A2(_02972_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08716_ (.A1(_02452_),
    .A2(_02974_),
    .B(_02979_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08717_ (.A1(_02402_),
    .A2(_02970_),
    .B1(_02983_),
    .B2(_02984_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08718_ (.I(_02710_),
    .Z(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08719_ (.A1(\as2650.stack[15][4] ),
    .A2(_02972_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08720_ (.A1(_02456_),
    .A2(_02712_),
    .B(_02979_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08721_ (.A1(_02405_),
    .A2(_02985_),
    .B1(_02986_),
    .B2(_02987_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08722_ (.A1(\as2650.stack[15][5] ),
    .A2(_02978_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08723_ (.I(_02109_),
    .Z(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08724_ (.A1(_02989_),
    .A2(_02712_),
    .B(_02969_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08725_ (.A1(_02409_),
    .A2(_02985_),
    .B1(_02988_),
    .B2(_02990_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08726_ (.A1(\as2650.stack[15][6] ),
    .A2(_02978_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08727_ (.A1(_02461_),
    .A2(_02712_),
    .B(_02969_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08728_ (.A1(_02412_),
    .A2(_02985_),
    .B1(_02991_),
    .B2(_02992_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08729_ (.A1(_02381_),
    .A2(_02974_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08730_ (.A1(\as2650.stack[15][7] ),
    .A2(_02978_),
    .B(_02969_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08731_ (.A1(_02415_),
    .A2(_02985_),
    .B1(_02993_),
    .B2(_02994_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08732_ (.I(_02692_),
    .Z(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08733_ (.I(_02995_),
    .Z(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08734_ (.A1(_02003_),
    .A2(_02437_),
    .A3(_02147_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08735_ (.I(_02997_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08736_ (.A1(\as2650.stack[1][0] ),
    .A2(_02998_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08737_ (.I(_02044_),
    .Z(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08738_ (.I(_02688_),
    .Z(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08739_ (.A1(_03000_),
    .A2(_03001_),
    .B(_02701_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08740_ (.A1(_02384_),
    .A2(_02996_),
    .B1(_02999_),
    .B2(_03002_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08741_ (.A1(_02976_),
    .A2(_02700_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08742_ (.I(_02997_),
    .Z(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08743_ (.I(_02693_),
    .Z(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08744_ (.A1(\as2650.stack[1][1] ),
    .A2(_03004_),
    .B(_03005_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08745_ (.A1(_02394_),
    .A2(_02996_),
    .B1(_03003_),
    .B2(_03006_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08746_ (.A1(\as2650.stack[1][2] ),
    .A2(_02998_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08747_ (.A1(_02449_),
    .A2(_03001_),
    .B(_03005_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08748_ (.A1(_02399_),
    .A2(_02996_),
    .B1(_03007_),
    .B2(_03008_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08749_ (.A1(\as2650.stack[1][3] ),
    .A2(_02998_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08750_ (.A1(_02452_),
    .A2(_03001_),
    .B(_03005_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08751_ (.A1(_02402_),
    .A2(_02996_),
    .B1(_03009_),
    .B2(_03010_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08752_ (.I(_02693_),
    .Z(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08753_ (.A1(_02097_),
    .A2(_03001_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08754_ (.A1(\as2650.stack[1][4] ),
    .A2(_03004_),
    .B(_03005_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08755_ (.A1(_02405_),
    .A2(_03011_),
    .B1(_03012_),
    .B2(_03013_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08756_ (.A1(\as2650.stack[1][5] ),
    .A2(_02998_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08757_ (.A1(_02989_),
    .A2(_02695_),
    .B(_02995_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08758_ (.A1(_02409_),
    .A2(_03011_),
    .B1(_03014_),
    .B2(_03015_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08759_ (.A1(\as2650.stack[1][6] ),
    .A2(_03004_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08760_ (.A1(_02461_),
    .A2(_02695_),
    .B(_02995_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08761_ (.A1(_02412_),
    .A2(_03011_),
    .B1(_03016_),
    .B2(_03017_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08762_ (.A1(\as2650.stack[1][7] ),
    .A2(_03004_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08763_ (.A1(_02302_),
    .A2(_02695_),
    .B(_02995_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08764_ (.A1(_02415_),
    .A2(_03011_),
    .B1(_03018_),
    .B2(_03019_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08765_ (.I(_01983_),
    .Z(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08766_ (.I(_02472_),
    .Z(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08767_ (.I(_03021_),
    .Z(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08768_ (.A1(_02151_),
    .A2(_02480_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08769_ (.I(_02022_),
    .Z(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08770_ (.A1(_02388_),
    .A2(_02146_),
    .A3(_03024_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08771_ (.I(_03025_),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08772_ (.A1(\as2650.stack[8][0] ),
    .A2(_03026_),
    .B(_02481_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08773_ (.A1(_03020_),
    .A2(_03022_),
    .B1(_03023_),
    .B2(_03027_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08774_ (.I(_02050_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08775_ (.I(_02466_),
    .Z(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08776_ (.A1(_02976_),
    .A2(_03029_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08777_ (.I(_02473_),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08778_ (.A1(\as2650.stack[8][1] ),
    .A2(_03026_),
    .B(_03031_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08779_ (.A1(_03028_),
    .A2(_03022_),
    .B1(_03030_),
    .B2(_03032_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08780_ (.I(_02066_),
    .Z(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08781_ (.A1(_02368_),
    .A2(_03029_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08782_ (.I(_03025_),
    .Z(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08783_ (.A1(\as2650.stack[8][2] ),
    .A2(_03035_),
    .B(_03031_),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08784_ (.A1(_03033_),
    .A2(_03022_),
    .B1(_03034_),
    .B2(_03036_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08785_ (.I(_02077_),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08786_ (.A1(\as2650.stack[8][3] ),
    .A2(_03026_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08787_ (.A1(_02452_),
    .A2(_02475_),
    .B(_03031_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08788_ (.A1(_03037_),
    .A2(_03022_),
    .B1(_03038_),
    .B2(_03039_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08789_ (.I(_02090_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08790_ (.I(_02473_),
    .Z(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08791_ (.A1(_02097_),
    .A2(_03029_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08792_ (.A1(\as2650.stack[8][4] ),
    .A2(_03035_),
    .B(_03031_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08793_ (.A1(_03040_),
    .A2(_03041_),
    .B1(_03042_),
    .B2(_03043_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08794_ (.I(_02101_),
    .Z(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08795_ (.A1(_02376_),
    .A2(_03029_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08796_ (.A1(\as2650.stack[8][5] ),
    .A2(_03035_),
    .B(_03021_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08797_ (.A1(_03044_),
    .A2(_03041_),
    .B1(_03045_),
    .B2(_03046_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08798_ (.I(_02112_),
    .Z(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08799_ (.A1(\as2650.stack[8][6] ),
    .A2(_03026_),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08800_ (.A1(_02461_),
    .A2(_02475_),
    .B(_03021_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08801_ (.A1(_03047_),
    .A2(_03041_),
    .B1(_03048_),
    .B2(_03049_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08802_ (.I(_02121_),
    .Z(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08803_ (.A1(_02381_),
    .A2(_02475_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08804_ (.A1(\as2650.stack[8][7] ),
    .A2(_03035_),
    .B(_03021_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08805_ (.A1(_03050_),
    .A2(_03041_),
    .B1(_03051_),
    .B2(_03052_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08806_ (.A1(_00940_),
    .A2(_00651_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08807_ (.I(_03053_),
    .Z(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08808_ (.A1(_00945_),
    .A2(_03054_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08809_ (.A1(_01050_),
    .A2(_03054_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08810_ (.I(_03056_),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08811_ (.A1(_00923_),
    .A2(_00927_),
    .A3(_00931_),
    .A4(_03053_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08812_ (.I(_03058_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08813_ (.A1(_00953_),
    .A2(_03055_),
    .B(_03057_),
    .C(_03059_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08814_ (.A1(_00955_),
    .A2(_00941_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08815_ (.A1(_01129_),
    .A2(_01131_),
    .A3(_03061_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08816_ (.I(_03062_),
    .Z(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08817_ (.A1(_02089_),
    .A2(_00982_),
    .A3(_00967_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08818_ (.I(_03064_),
    .Z(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08819_ (.A1(_00987_),
    .A2(_00995_),
    .A3(_03054_),
    .Z(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08820_ (.A1(_03060_),
    .A2(_03063_),
    .A3(_03065_),
    .A4(_03066_),
    .Z(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08821_ (.A1(_00921_),
    .A2(_03067_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08822_ (.I(_03065_),
    .Z(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08823_ (.I(_03066_),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08824_ (.I(_03070_),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08825_ (.A1(_00981_),
    .A2(_00983_),
    .A3(_03054_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08826_ (.I(_03072_),
    .Z(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08827_ (.I(_03072_),
    .Z(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08828_ (.I(_03057_),
    .Z(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08829_ (.A1(_00744_),
    .A2(_00937_),
    .A3(_03061_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08830_ (.A1(_01026_),
    .A2(_03076_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08831_ (.I(_03077_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08832_ (.A1(_01143_),
    .A2(_03076_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08833_ (.I(_03079_),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08834_ (.A1(_01604_),
    .A2(_03061_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08835_ (.I(_03081_),
    .Z(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08836_ (.A1(_01043_),
    .A2(_03082_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08837_ (.A1(_00428_),
    .A2(_03082_),
    .B(_03079_),
    .C(_03083_),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08838_ (.I(_03077_),
    .Z(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08839_ (.A1(_01277_),
    .A2(_03080_),
    .B(_03084_),
    .C(_03085_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08840_ (.I(_03056_),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08841_ (.A1(_01032_),
    .A2(_03078_),
    .B(_03086_),
    .C(_03087_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08842_ (.A1(_01100_),
    .A2(_03075_),
    .B(_03088_),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08843_ (.A1(_03074_),
    .A2(_03089_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08844_ (.A1(_01019_),
    .A2(_03073_),
    .B(_03090_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08845_ (.A1(_01120_),
    .A2(_01010_),
    .Z(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08846_ (.I(_03070_),
    .Z(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08847_ (.A1(_03092_),
    .A2(_03093_),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08848_ (.A1(_03071_),
    .A2(_03091_),
    .B(_03094_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08849_ (.I(_03065_),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08850_ (.A1(_01097_),
    .A2(_03096_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08851_ (.A1(_03069_),
    .A2(_03095_),
    .B(_03097_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08852_ (.A1(_00921_),
    .A2(_03067_),
    .Z(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08853_ (.A1(_00606_),
    .A2(_00745_),
    .A3(_01024_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08854_ (.A1(_01103_),
    .A2(_03100_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08855_ (.A1(_00835_),
    .A2(_03101_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08856_ (.I(_03102_),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08857_ (.A1(_00695_),
    .A2(_03099_),
    .A3(_03103_),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08858_ (.I(_03104_),
    .Z(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08859_ (.A1(\as2650.r123_2[1][0] ),
    .A2(_03105_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08860_ (.I(_03103_),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08861_ (.I(_03107_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08862_ (.A1(_01102_),
    .A2(_01112_),
    .A3(_03108_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08863_ (.A1(_03068_),
    .A2(_03098_),
    .B(_03106_),
    .C(_03109_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08864_ (.I(_03068_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08865_ (.I(_03057_),
    .Z(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08866_ (.I(_03077_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08867_ (.I(_03079_),
    .Z(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08868_ (.I(_03081_),
    .Z(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08869_ (.A1(_00609_),
    .A2(_03055_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08870_ (.A1(_01142_),
    .A2(_03082_),
    .B(_03115_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08871_ (.A1(_01146_),
    .A2(_03114_),
    .B(_03116_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08872_ (.A1(_01150_),
    .A2(_03113_),
    .B(_03117_),
    .C(_03085_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08873_ (.I(_03057_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08874_ (.A1(_01139_),
    .A2(_03112_),
    .B(_03118_),
    .C(_03119_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08875_ (.A1(_01136_),
    .A2(_03111_),
    .B(_03072_),
    .C(_03120_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08876_ (.I(_03062_),
    .Z(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08877_ (.A1(_01161_),
    .A2(_03122_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08878_ (.A1(_03121_),
    .A2(_03123_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08879_ (.I(_03070_),
    .Z(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08880_ (.I0(_03124_),
    .I1(_01127_),
    .S(_03125_),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08881_ (.I(_03065_),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08882_ (.A1(_01195_),
    .A2(_03127_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08883_ (.A1(_03069_),
    .A2(_03126_),
    .B(_03128_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08884_ (.I(_03104_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08885_ (.A1(_01206_),
    .A2(_03108_),
    .B1(_03130_),
    .B2(\as2650.r123_2[1][1] ),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08886_ (.A1(_03110_),
    .A2(_03129_),
    .B(_03131_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08887_ (.A1(_01262_),
    .A2(_03075_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08888_ (.I(_03077_),
    .Z(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08889_ (.I(_03059_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08890_ (.A1(_00426_),
    .A2(_03134_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08891_ (.A1(_02849_),
    .A2(_03059_),
    .B(_03113_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08892_ (.A1(_01297_),
    .A2(_03113_),
    .B1(_03135_),
    .B2(_03136_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08893_ (.I(_01034_),
    .Z(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08894_ (.A1(_03138_),
    .A2(_03112_),
    .B(_03087_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08895_ (.A1(_03133_),
    .A2(_03137_),
    .B(_03139_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08896_ (.A1(_01286_),
    .A2(_03063_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08897_ (.A1(_03122_),
    .A2(_03132_),
    .A3(_03140_),
    .B(_03141_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08898_ (.I0(_03142_),
    .I1(_01261_),
    .S(_03125_),
    .Z(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08899_ (.A1(_01249_),
    .A2(_03096_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08900_ (.A1(_03069_),
    .A2(_03143_),
    .B(_03144_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08901_ (.A1(_01222_),
    .A2(_03108_),
    .B1(_03130_),
    .B2(\as2650.r123_2[1][2] ),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08902_ (.A1(_03110_),
    .A2(_03145_),
    .B(_03146_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08903_ (.A1(_01156_),
    .A2(_01298_),
    .B1(_01300_),
    .B2(_01318_),
    .C(_01320_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08904_ (.I(_01234_),
    .Z(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08905_ (.I(_01309_),
    .Z(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08906_ (.I(_01310_),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08907_ (.I(_03058_),
    .Z(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08908_ (.A1(_00439_),
    .A2(_03058_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08909_ (.A1(_03150_),
    .A2(_03151_),
    .B(_03079_),
    .C(_03152_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08910_ (.A1(_03149_),
    .A2(_03080_),
    .B(_03153_),
    .C(_03085_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08911_ (.A1(_03148_),
    .A2(_03078_),
    .B(_03154_),
    .C(_03087_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08912_ (.A1(_01306_),
    .A2(_03075_),
    .B(_03155_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08913_ (.A1(_03074_),
    .A2(_03156_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08914_ (.A1(_03147_),
    .A2(_03073_),
    .B(_03157_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08915_ (.A1(_01303_),
    .A2(_03093_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08916_ (.A1(_03071_),
    .A2(_03158_),
    .B(_03159_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08917_ (.A1(_01350_),
    .A2(_03096_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08918_ (.A1(_03069_),
    .A2(_03160_),
    .B(_03161_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08919_ (.I(_03103_),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08920_ (.A1(_01370_),
    .A2(_03163_),
    .B1(_03130_),
    .B2(\as2650.r123_2[1][3] ),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08921_ (.A1(_03110_),
    .A2(_03162_),
    .B(_03164_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08922_ (.I(_01436_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08923_ (.A1(_05813_),
    .A2(_03151_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08924_ (.A1(_03165_),
    .A2(_03151_),
    .B(_03080_),
    .C(_03166_),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08925_ (.A1(_01599_),
    .A2(_03113_),
    .B(_03167_),
    .C(_03078_),
    .ZN(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08926_ (.A1(_01431_),
    .A2(_03133_),
    .B(_03168_),
    .C(_03119_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08927_ (.A1(_01430_),
    .A2(_03111_),
    .B(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08928_ (.A1(_01445_),
    .A2(_03074_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08929_ (.A1(_03073_),
    .A2(_03170_),
    .B(_03171_),
    .C(_03070_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08930_ (.A1(_01429_),
    .A2(_03093_),
    .B(_03172_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08931_ (.I0(_03173_),
    .I1(_01422_),
    .S(_03127_),
    .Z(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08932_ (.A1(_01387_),
    .A2(_03163_),
    .B1(_03130_),
    .B2(\as2650.r123_2[1][4] ),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08933_ (.A1(_03110_),
    .A2(_03174_),
    .B(_03175_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08934_ (.A1(\as2650.r123_2[1][5] ),
    .A2(_03105_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08935_ (.I(_03107_),
    .Z(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08936_ (.I(_03096_),
    .Z(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08937_ (.A1(_02836_),
    .A2(_03080_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08938_ (.A1(_05804_),
    .A2(_03082_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08939_ (.A1(_02933_),
    .A2(_03114_),
    .B(_03115_),
    .C(_03180_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08940_ (.A1(_03179_),
    .A2(_03181_),
    .B(_03085_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08941_ (.A1(_01460_),
    .A2(_03112_),
    .B(_03182_),
    .C(_03087_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08942_ (.A1(_01954_),
    .A2(_03111_),
    .B(_03072_),
    .C(_03183_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08943_ (.A1(_01474_),
    .A2(_03063_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08944_ (.A1(_03184_),
    .A2(_03185_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08945_ (.I0(_03186_),
    .I1(_01458_),
    .S(_03125_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08946_ (.A1(_03178_),
    .A2(_03187_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08947_ (.A1(_01501_),
    .A2(_03178_),
    .B(_03188_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08948_ (.A1(_01530_),
    .A2(_03177_),
    .B1(_03189_),
    .B2(_03099_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08949_ (.A1(_03176_),
    .A2(_03190_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08950_ (.A1(\as2650.r123_2[1][6] ),
    .A2(_03105_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08951_ (.I(_03115_),
    .Z(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08952_ (.A1(_05801_),
    .A2(_03059_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08953_ (.A1(_01611_),
    .A2(_03114_),
    .B(_03192_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08954_ (.A1(_01602_),
    .A2(_03192_),
    .B1(_03193_),
    .B2(_03194_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08955_ (.A1(_03112_),
    .A2(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08956_ (.A1(_02835_),
    .A2(_03133_),
    .B(_03196_),
    .C(_03075_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08957_ (.A1(_01597_),
    .A2(_03119_),
    .Z(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08958_ (.A1(_03197_),
    .A2(_03198_),
    .B(_03122_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08959_ (.A1(_01596_),
    .A2(_03122_),
    .B(_03125_),
    .C(_03199_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08960_ (.A1(_01619_),
    .A2(_03071_),
    .B(_03200_),
    .C(_03127_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08961_ (.A1(_01589_),
    .A2(_03178_),
    .B(_03201_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08962_ (.A1(_01563_),
    .A2(_03177_),
    .B1(_03202_),
    .B2(_03099_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08963_ (.A1(_03191_),
    .A2(_03203_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08964_ (.A1(\as2650.r123_2[1][7] ),
    .A2(_03105_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08965_ (.A1(_05796_),
    .A2(_03151_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08966_ (.A1(_02932_),
    .A2(_03114_),
    .B(_03192_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08967_ (.A1(_01700_),
    .A2(_03192_),
    .B1(_03205_),
    .B2(_03206_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08968_ (.A1(_03078_),
    .A2(_03207_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08969_ (.A1(_02836_),
    .A2(_03133_),
    .B(_03208_),
    .C(_03119_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08970_ (.A1(_02345_),
    .A2(_03111_),
    .B(_03209_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08971_ (.A1(_01696_),
    .A2(_03074_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08972_ (.A1(_03073_),
    .A2(_03210_),
    .B(_03211_),
    .C(_03093_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08973_ (.A1(_01693_),
    .A2(_03071_),
    .B(_03212_),
    .C(_03127_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08974_ (.A1(_01686_),
    .A2(_03178_),
    .B(_03213_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08975_ (.A1(_01658_),
    .A2(_03177_),
    .B1(_03214_),
    .B2(_03099_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08976_ (.A1(_03204_),
    .A2(_03215_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08977_ (.I(_02492_),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08978_ (.I(_03216_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08979_ (.A1(_02648_),
    .A2(_02000_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08980_ (.A1(_02143_),
    .A2(_02438_),
    .A3(_03218_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08981_ (.I(_03219_),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08982_ (.A1(\as2650.stack[7][0] ),
    .A2(_03220_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08983_ (.I(_02487_),
    .Z(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08984_ (.A1(_03000_),
    .A2(_03222_),
    .B(_02501_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08985_ (.A1(_03020_),
    .A2(_03217_),
    .B1(_03221_),
    .B2(_03223_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08986_ (.A1(\as2650.stack[7][1] ),
    .A2(_03220_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08987_ (.I(_02493_),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08988_ (.A1(_02364_),
    .A2(_03222_),
    .B(_03225_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08989_ (.A1(_03028_),
    .A2(_03217_),
    .B1(_03224_),
    .B2(_03226_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08990_ (.A1(_02368_),
    .A2(_02500_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08991_ (.I(_03219_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08992_ (.A1(\as2650.stack[7][2] ),
    .A2(_03228_),
    .B(_03225_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08993_ (.A1(_03033_),
    .A2(_03217_),
    .B1(_03227_),
    .B2(_03229_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08994_ (.A1(\as2650.stack[7][3] ),
    .A2(_03220_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08995_ (.I(_02086_),
    .Z(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08996_ (.A1(_03231_),
    .A2(_03222_),
    .B(_03225_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08997_ (.A1(_03037_),
    .A2(_03217_),
    .B1(_03230_),
    .B2(_03232_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08998_ (.I(_02493_),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08999_ (.A1(_02097_),
    .A2(_03222_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09000_ (.A1(\as2650.stack[7][4] ),
    .A2(_03228_),
    .B(_03225_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09001_ (.A1(_03040_),
    .A2(_03233_),
    .B1(_03234_),
    .B2(_03235_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09002_ (.A1(\as2650.stack[7][5] ),
    .A2(_03220_),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09003_ (.A1(_02989_),
    .A2(_02495_),
    .B(_03216_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09004_ (.A1(_03044_),
    .A2(_03233_),
    .B1(_03236_),
    .B2(_03237_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09005_ (.A1(\as2650.stack[7][6] ),
    .A2(_03228_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09006_ (.I(_02118_),
    .Z(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09007_ (.A1(_03239_),
    .A2(_02495_),
    .B(_03216_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09008_ (.A1(_03047_),
    .A2(_03233_),
    .B1(_03238_),
    .B2(_03240_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09009_ (.A1(\as2650.stack[7][7] ),
    .A2(_03228_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09010_ (.A1(_02302_),
    .A2(_02495_),
    .B(_03216_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09011_ (.A1(_03050_),
    .A2(_03233_),
    .B1(_03241_),
    .B2(_03242_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09012_ (.A1(_05696_),
    .A2(_00826_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09013_ (.A1(_03243_),
    .A2(_03067_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09014_ (.I(_03244_),
    .Z(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09015_ (.A1(_00848_),
    .A2(_03101_),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09016_ (.A1(_03102_),
    .A2(_03246_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09017_ (.I(_03247_),
    .Z(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09018_ (.A1(_01725_),
    .A2(_03101_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09019_ (.I(_03249_),
    .Z(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09020_ (.I(_03250_),
    .Z(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09021_ (.I(_03249_),
    .Z(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09022_ (.A1(_01800_),
    .A2(_03252_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09023_ (.A1(_01101_),
    .A2(_03251_),
    .B(_03253_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09024_ (.A1(_03098_),
    .A2(_03245_),
    .B1(_03248_),
    .B2(_03254_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09025_ (.A1(_03060_),
    .A2(_03063_),
    .A3(_03064_),
    .A4(_03066_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09026_ (.A1(_00838_),
    .A2(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09027_ (.A1(_05677_),
    .A2(_03257_),
    .A3(_03246_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09028_ (.I(_03258_),
    .Z(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09029_ (.I0(_03255_),
    .I1(\as2650.r123_2[0][0] ),
    .S(_03259_),
    .Z(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09030_ (.I(_03260_),
    .Z(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09031_ (.I(_01203_),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09032_ (.I(_03249_),
    .Z(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09033_ (.A1(_01847_),
    .A2(_03252_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09034_ (.A1(_03261_),
    .A2(_03262_),
    .B(_03263_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09035_ (.A1(_03129_),
    .A2(_03245_),
    .B1(_03248_),
    .B2(_03264_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09036_ (.I0(_03265_),
    .I1(\as2650.r123_2[0][1] ),
    .S(_03259_),
    .Z(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09037_ (.I(_03266_),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09038_ (.I(_01263_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09039_ (.A1(_01884_),
    .A2(_03250_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09040_ (.A1(_03267_),
    .A2(_03262_),
    .B(_03268_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09041_ (.A1(_03145_),
    .A2(_03245_),
    .B1(_03248_),
    .B2(_03269_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09042_ (.I(_03258_),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09043_ (.I0(_03270_),
    .I1(\as2650.r123_2[0][2] ),
    .S(_03271_),
    .Z(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09044_ (.I(_03272_),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09045_ (.I(_01905_),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09046_ (.A1(_01904_),
    .A2(_03250_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09047_ (.A1(_03273_),
    .A2(_03262_),
    .B(_03274_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09048_ (.A1(_03162_),
    .A2(_03245_),
    .B1(_03248_),
    .B2(_03275_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09049_ (.I0(_03276_),
    .I1(\as2650.r123_2[0][3] ),
    .S(_03271_),
    .Z(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09050_ (.I(_03277_),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09051_ (.I(_03247_),
    .Z(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09052_ (.I(_01927_),
    .Z(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09053_ (.A1(_01926_),
    .A2(_03250_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09054_ (.A1(_03279_),
    .A2(_03262_),
    .B(_03280_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09055_ (.A1(_03174_),
    .A2(_03244_),
    .B1(_03278_),
    .B2(_03281_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09056_ (.I0(_03282_),
    .I1(\as2650.r123_2[0][4] ),
    .S(_03271_),
    .Z(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09057_ (.I(_03283_),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09058_ (.I(_03271_),
    .Z(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09059_ (.I(_01954_),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09060_ (.A1(_03285_),
    .A2(_03252_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09061_ (.A1(_01953_),
    .A2(_03251_),
    .B(_03278_),
    .C(_03286_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09062_ (.A1(_03189_),
    .A2(_03257_),
    .B(_03287_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09063_ (.A1(\as2650.r123_2[0][5] ),
    .A2(_03284_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09064_ (.A1(_03284_),
    .A2(_03288_),
    .B(_03289_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09065_ (.A1(_01975_),
    .A2(_03252_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09066_ (.A1(_01974_),
    .A2(_03251_),
    .B(_03278_),
    .C(_03290_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09067_ (.A1(_03202_),
    .A2(_03257_),
    .B(_03291_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09068_ (.A1(\as2650.r123_2[0][6] ),
    .A2(_03259_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09069_ (.A1(_03284_),
    .A2(_03292_),
    .B(_03293_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09070_ (.A1(_01980_),
    .A2(_03251_),
    .A3(_03278_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09071_ (.A1(_03214_),
    .A2(_03257_),
    .B(_03294_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09072_ (.A1(\as2650.r123_2[0][7] ),
    .A2(_03259_),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09073_ (.A1(_03284_),
    .A2(_03295_),
    .B(_03296_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09074_ (.A1(_00514_),
    .A2(_03067_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09075_ (.I(_03297_),
    .Z(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09076_ (.A1(_01628_),
    .A2(_01656_),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09077_ (.A1(_01626_),
    .A2(_01657_),
    .B(_03299_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09078_ (.A1(_01634_),
    .A2(_01654_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09079_ (.A1(_01631_),
    .A2(_01655_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09080_ (.A1(_03301_),
    .A2(_03302_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09081_ (.A1(_01569_),
    .A2(_01204_),
    .A3(_01637_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09082_ (.A1(_01639_),
    .A2(_01640_),
    .B(_03304_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09083_ (.A1(_01547_),
    .A2(_01551_),
    .A3(_01652_),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09084_ (.A1(_01641_),
    .A2(_01653_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09085_ (.A1(_03306_),
    .A2(_03307_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09086_ (.A1(_01635_),
    .A2(_01644_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09087_ (.A1(_05758_),
    .A2(_01379_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09088_ (.A1(_01550_),
    .A2(_03310_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09089_ (.A1(_01643_),
    .A2(_03309_),
    .B(_03311_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09090_ (.A1(_05723_),
    .A2(_01212_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09091_ (.A1(_03312_),
    .A2(_03313_),
    .Z(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09092_ (.A1(_03312_),
    .A2(_03313_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09093_ (.A1(_03314_),
    .A2(_03315_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09094_ (.A1(_01546_),
    .A2(_01651_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09095_ (.A1(_01546_),
    .A2(_01651_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09096_ (.A1(_01645_),
    .A2(_03317_),
    .B(_03318_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09097_ (.A1(\as2650.r0[1] ),
    .A2(_01648_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09098_ (.A1(_05780_),
    .A2(_01543_),
    .B1(_01649_),
    .B2(\as2650.r0[0] ),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09099_ (.A1(_01544_),
    .A2(_03320_),
    .B1(_03321_),
    .B2(_01647_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09100_ (.A1(\as2650.r0[2] ),
    .A2(_01542_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09101_ (.A1(_05764_),
    .A2(_01515_),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09102_ (.A1(_03320_),
    .A2(_03323_),
    .A3(_03324_),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09103_ (.A1(_03322_),
    .A2(_03325_),
    .Z(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09104_ (.A1(\as2650.r0[6] ),
    .A2(_01217_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09105_ (.A1(_05731_),
    .A2(_01358_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09106_ (.A1(_03310_),
    .A2(_03328_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09107_ (.A1(_03327_),
    .A2(_03329_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09108_ (.A1(_03326_),
    .A2(_03330_),
    .Z(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09109_ (.A1(_03319_),
    .A2(_03331_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09110_ (.A1(_03316_),
    .A2(_03332_),
    .Z(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09111_ (.A1(_03308_),
    .A2(_03333_),
    .Z(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09112_ (.A1(_03305_),
    .A2(_03334_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09113_ (.A1(_03303_),
    .A2(_03335_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09114_ (.A1(_03300_),
    .A2(_03336_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09115_ (.A1(_05697_),
    .A2(_03256_),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09116_ (.A1(_00640_),
    .A2(_03103_),
    .A3(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09117_ (.I(_03339_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09118_ (.A1(_03108_),
    .A2(_03337_),
    .B1(_03340_),
    .B2(\as2650.r123_2[2][0] ),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09119_ (.A1(_03098_),
    .A2(_03298_),
    .B(_03341_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09120_ (.I(_03339_),
    .Z(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09121_ (.A1(_03303_),
    .A2(_03335_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09122_ (.A1(_03300_),
    .A2(_03336_),
    .B(_03343_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09123_ (.A1(_03308_),
    .A2(_03333_),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09124_ (.A1(_03305_),
    .A2(_03334_),
    .B(_03345_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09125_ (.A1(_03319_),
    .A2(_03331_),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09126_ (.A1(_03316_),
    .A2(_03332_),
    .B(_03347_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09127_ (.A1(_05731_),
    .A2(_01510_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09128_ (.A1(_01644_),
    .A2(_03349_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09129_ (.A1(_03327_),
    .A2(_03329_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09130_ (.A1(_03350_),
    .A2(_03351_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09131_ (.I(_03322_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09132_ (.A1(_03326_),
    .A2(_03330_),
    .Z(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09133_ (.A1(_03353_),
    .A2(_03325_),
    .B(_03354_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09134_ (.A1(_03320_),
    .A2(_03323_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09135_ (.A1(_05750_),
    .A2(_01649_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09136_ (.A1(_01646_),
    .A2(_03357_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09137_ (.A1(_03356_),
    .A2(_03324_),
    .B(_03358_),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09138_ (.A1(_05764_),
    .A2(_01542_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09139_ (.A1(_03357_),
    .A2(_03360_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09140_ (.A1(_05759_),
    .A2(_01516_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09141_ (.A1(_03361_),
    .A2(_03362_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09142_ (.A1(_03359_),
    .A2(_03363_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09143_ (.A1(\as2650.r0[7] ),
    .A2(_01218_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09144_ (.A1(_05742_),
    .A2(_01360_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09145_ (.A1(_03349_),
    .A2(_03366_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09146_ (.A1(_03365_),
    .A2(_03367_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09147_ (.A1(_03364_),
    .A2(_03368_),
    .Z(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09148_ (.A1(_03355_),
    .A2(_03369_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09149_ (.A1(_03352_),
    .A2(_03370_),
    .Z(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09150_ (.A1(_03314_),
    .A2(_03348_),
    .A3(_03371_),
    .Z(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09151_ (.A1(_03346_),
    .A2(_03372_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09152_ (.A1(_03344_),
    .A2(_03373_),
    .Z(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09153_ (.A1(\as2650.r123_2[2][1] ),
    .A2(_03342_),
    .B1(_03374_),
    .B2(_03163_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09154_ (.A1(_03129_),
    .A2(_03298_),
    .B(_03375_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09155_ (.A1(_03346_),
    .A2(_03372_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09156_ (.A1(_03344_),
    .A2(_03373_),
    .B(_03376_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09157_ (.A1(_03348_),
    .A2(_03371_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09158_ (.A1(_03348_),
    .A2(_03371_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09159_ (.A1(_03314_),
    .A2(_03378_),
    .B(_03379_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09160_ (.A1(_03355_),
    .A2(_03369_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09161_ (.A1(_03352_),
    .A2(_03370_),
    .B(_03381_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09162_ (.A1(_03349_),
    .A2(_03366_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09163_ (.A1(_03365_),
    .A2(_03367_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09164_ (.A1(_03383_),
    .A2(_03384_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09165_ (.A1(_03364_),
    .A2(_03368_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09166_ (.A1(_03359_),
    .A2(_03363_),
    .B(_03386_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09167_ (.A1(_05724_),
    .A2(_01363_),
    .B1(_02223_),
    .B2(_05743_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09168_ (.A1(_05723_),
    .A2(_01380_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09169_ (.A1(_03366_),
    .A2(_03389_),
    .Z(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09170_ (.I(_03390_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09171_ (.A1(_03388_),
    .A2(_03391_),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09172_ (.I(_01649_),
    .Z(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09173_ (.A1(_05765_),
    .A2(_03393_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09174_ (.A1(_03323_),
    .A2(_03394_),
    .B1(_03361_),
    .B2(_03362_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09175_ (.A1(_05758_),
    .A2(_02233_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09176_ (.A1(_03394_),
    .A2(_03396_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09177_ (.A1(_05732_),
    .A2(_01517_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09178_ (.A1(_03397_),
    .A2(_03398_),
    .Z(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09179_ (.A1(_03395_),
    .A2(_03399_),
    .Z(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09180_ (.A1(_03392_),
    .A2(_03400_),
    .Z(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09181_ (.A1(_03387_),
    .A2(_03401_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09182_ (.A1(_03385_),
    .A2(_03402_),
    .Z(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09183_ (.A1(_03382_),
    .A2(_03403_),
    .Z(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09184_ (.A1(_03380_),
    .A2(_03404_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09185_ (.A1(_03377_),
    .A2(_03405_),
    .Z(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09186_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_03342_),
    .B1(_03406_),
    .B2(_03163_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09187_ (.A1(_03145_),
    .A2(_03298_),
    .B(_03407_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09188_ (.A1(_03380_),
    .A2(_03404_),
    .Z(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09189_ (.A1(_03377_),
    .A2(_03405_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09190_ (.A1(_03408_),
    .A2(_03409_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09191_ (.A1(_03382_),
    .A2(_03403_),
    .Z(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09192_ (.A1(_03395_),
    .A2(_03399_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09193_ (.A1(_03392_),
    .A2(_03400_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09194_ (.A1(_03412_),
    .A2(_03413_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09195_ (.A1(_05759_),
    .A2(_03393_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09196_ (.A1(_03360_),
    .A2(_03415_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09197_ (.A1(_03397_),
    .A2(_03398_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09198_ (.A1(_03416_),
    .A2(_03417_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09199_ (.A1(_05731_),
    .A2(_02233_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09200_ (.A1(_03415_),
    .A2(_03419_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09201_ (.A1(_05743_),
    .A2(_01517_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09202_ (.A1(_03420_),
    .A2(_03421_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09203_ (.A1(_03418_),
    .A2(_03422_),
    .Z(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09204_ (.A1(_03389_),
    .A2(_03423_),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09205_ (.A1(_03414_),
    .A2(_03424_),
    .Z(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09206_ (.A1(_03390_),
    .A2(_03425_),
    .Z(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09207_ (.A1(_03387_),
    .A2(_03401_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09208_ (.A1(_03385_),
    .A2(_03402_),
    .B(_03427_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09209_ (.A1(_03426_),
    .A2(_03428_),
    .Z(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09210_ (.A1(_03411_),
    .A2(_03429_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09211_ (.A1(_03410_),
    .A2(_03430_),
    .Z(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09212_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_03342_),
    .B1(_03431_),
    .B2(_03107_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09213_ (.A1(_03162_),
    .A2(_03298_),
    .B(_03432_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09214_ (.A1(_03411_),
    .A2(_03408_),
    .B(_03429_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09215_ (.A1(_03377_),
    .A2(_03405_),
    .A3(_03430_),
    .B(_03433_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09216_ (.A1(_03426_),
    .A2(_03428_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09217_ (.A1(_05733_),
    .A2(_03393_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09218_ (.A1(_03396_),
    .A2(_03436_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09219_ (.A1(_03420_),
    .A2(_03421_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09220_ (.A1(_03437_),
    .A2(_03438_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09221_ (.A1(_01569_),
    .A2(_02233_),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09222_ (.A1(_03436_),
    .A2(_03440_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09223_ (.A1(_05724_),
    .A2(_01518_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09224_ (.A1(_03441_),
    .A2(_03442_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09225_ (.A1(_03439_),
    .A2(_03443_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09226_ (.A1(_01663_),
    .A2(_02223_),
    .A3(_03423_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09227_ (.A1(_03418_),
    .A2(_03422_),
    .B(_03445_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09228_ (.A1(_03444_),
    .A2(_03446_),
    .Z(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09229_ (.I(_03424_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09230_ (.A1(_03414_),
    .A2(_03448_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09231_ (.A1(_03390_),
    .A2(_03425_),
    .Z(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09232_ (.A1(_03449_),
    .A2(_03450_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09233_ (.A1(_03447_),
    .A2(_03451_),
    .Z(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09234_ (.A1(_03435_),
    .A2(_03452_),
    .Z(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09235_ (.A1(_03434_),
    .A2(_03453_),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09236_ (.A1(\as2650.r123_2[2][4] ),
    .A2(_03340_),
    .B1(_03454_),
    .B2(_03107_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09237_ (.A1(_03174_),
    .A2(_03297_),
    .B(_03455_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09238_ (.A1(_03189_),
    .A2(_03338_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09239_ (.A1(_03435_),
    .A2(_03452_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09240_ (.A1(_03435_),
    .A2(_03452_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09241_ (.A1(_03434_),
    .A2(_03457_),
    .B(_03458_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09242_ (.A1(_03449_),
    .A2(_03450_),
    .B(_03447_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09243_ (.A1(_03439_),
    .A2(_03443_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09244_ (.I(_03446_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09245_ (.A1(_03444_),
    .A2(_03462_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09246_ (.A1(_03461_),
    .A2(_03463_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09247_ (.I(_03393_),
    .Z(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09248_ (.A1(_01597_),
    .A2(_03465_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09249_ (.A1(_03419_),
    .A2(_03466_),
    .B1(_03441_),
    .B2(_03442_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09250_ (.A1(_01663_),
    .A2(_02234_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09251_ (.A1(_03466_),
    .A2(_03468_),
    .Z(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09252_ (.A1(_03467_),
    .A2(_03469_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09253_ (.A1(_03464_),
    .A2(_03470_),
    .Z(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09254_ (.A1(_03460_),
    .A2(_03471_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09255_ (.A1(_03459_),
    .A2(_03472_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09256_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_03342_),
    .B1(_03473_),
    .B2(_03177_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09257_ (.A1(_03456_),
    .A2(_03474_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09258_ (.A1(_00835_),
    .A2(_03101_),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09259_ (.A1(_03460_),
    .A2(_03471_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09260_ (.A1(_03459_),
    .A2(_03472_),
    .B(_03476_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09261_ (.I(_03470_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09262_ (.A1(_03463_),
    .A2(_03478_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09263_ (.A1(_02345_),
    .A2(_03465_),
    .A3(_03440_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09264_ (.A1(_03467_),
    .A2(_03469_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09265_ (.A1(_03439_),
    .A2(_03443_),
    .A3(_03470_),
    .B(_03481_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09266_ (.A1(_03480_),
    .A2(_03482_),
    .Z(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09267_ (.A1(_03477_),
    .A2(_03479_),
    .A3(_03483_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09268_ (.A1(_03202_),
    .A2(_03338_),
    .B1(_03340_),
    .B2(\as2650.r123_2[2][6] ),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09269_ (.A1(_03475_),
    .A2(_03484_),
    .B(_03485_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09270_ (.A1(_03479_),
    .A2(_03483_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09271_ (.A1(_02346_),
    .A2(_03465_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09272_ (.A1(_01975_),
    .A2(_02234_),
    .B(_03482_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09273_ (.A1(_03487_),
    .A2(_03488_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09274_ (.A1(_03479_),
    .A2(_03483_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09275_ (.A1(_03477_),
    .A2(_03486_),
    .B(_03489_),
    .C(_03490_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09276_ (.A1(_03214_),
    .A2(_03338_),
    .B1(_03340_),
    .B2(\as2650.r123_2[2][7] ),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09277_ (.A1(_03475_),
    .A2(_03491_),
    .B(_03492_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09278_ (.I(_02669_),
    .Z(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09279_ (.I(_03493_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09280_ (.A1(_02272_),
    .A2(_02437_),
    .A3(_03024_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09281_ (.I(_03495_),
    .Z(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09282_ (.A1(\as2650.stack[2][0] ),
    .A2(_03496_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09283_ (.A1(_03000_),
    .A2(_02673_),
    .B(_02682_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09284_ (.A1(_03020_),
    .A2(_03494_),
    .B1(_03497_),
    .B2(_03498_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09285_ (.A1(_02976_),
    .A2(_02681_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09286_ (.I(_02670_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09287_ (.A1(\as2650.stack[2][1] ),
    .A2(_03496_),
    .B(_03500_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09288_ (.A1(_03028_),
    .A2(_03494_),
    .B1(_03499_),
    .B2(_03501_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09289_ (.I(_02665_),
    .Z(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09290_ (.A1(_02368_),
    .A2(_03502_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09291_ (.I(_03495_),
    .Z(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09292_ (.A1(\as2650.stack[2][2] ),
    .A2(_03504_),
    .B(_03500_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09293_ (.A1(_03033_),
    .A2(_03494_),
    .B1(_03503_),
    .B2(_03505_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09294_ (.A1(\as2650.stack[2][3] ),
    .A2(_03496_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09295_ (.A1(_03231_),
    .A2(_02673_),
    .B(_03500_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09296_ (.A1(_03037_),
    .A2(_03494_),
    .B1(_03506_),
    .B2(_03507_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09297_ (.I(_02670_),
    .Z(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09298_ (.I(_02096_),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09299_ (.A1(_03509_),
    .A2(_03502_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09300_ (.A1(\as2650.stack[2][4] ),
    .A2(_03504_),
    .B(_03500_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09301_ (.A1(_03040_),
    .A2(_03508_),
    .B1(_03510_),
    .B2(_03511_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09302_ (.A1(_02376_),
    .A2(_03502_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09303_ (.A1(\as2650.stack[2][5] ),
    .A2(_03504_),
    .B(_03493_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09304_ (.A1(_03044_),
    .A2(_03508_),
    .B1(_03512_),
    .B2(_03513_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09305_ (.A1(\as2650.stack[2][6] ),
    .A2(_03496_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09306_ (.A1(_03239_),
    .A2(_02673_),
    .B(_03493_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09307_ (.A1(_03047_),
    .A2(_03508_),
    .B1(_03514_),
    .B2(_03515_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09308_ (.A1(_02184_),
    .A2(_03502_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09309_ (.A1(\as2650.stack[2][7] ),
    .A2(_03504_),
    .B(_03493_),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09310_ (.A1(_03050_),
    .A2(_03508_),
    .B1(_03516_),
    .B2(_03517_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09311_ (.I(_02631_),
    .Z(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09312_ (.I(_03518_),
    .Z(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09313_ (.A1(_02388_),
    .A2(_02438_),
    .A3(_03218_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09314_ (.I(_03520_),
    .Z(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09315_ (.A1(\as2650.stack[4][0] ),
    .A2(_03521_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09316_ (.I(_02626_),
    .Z(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09317_ (.A1(_03000_),
    .A2(_03523_),
    .B(_02640_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09318_ (.A1(_03020_),
    .A2(_03519_),
    .B1(_03522_),
    .B2(_03524_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09319_ (.A1(_02284_),
    .A2(_02639_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09320_ (.I(_03520_),
    .Z(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09321_ (.I(_02632_),
    .Z(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09322_ (.A1(\as2650.stack[4][1] ),
    .A2(_03526_),
    .B(_03527_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09323_ (.A1(_03028_),
    .A2(_03519_),
    .B1(_03525_),
    .B2(_03528_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09324_ (.A1(\as2650.stack[4][2] ),
    .A2(_03521_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09325_ (.A1(_02449_),
    .A2(_03523_),
    .B(_03527_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09326_ (.A1(_03033_),
    .A2(_03519_),
    .B1(_03529_),
    .B2(_03530_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09327_ (.A1(\as2650.stack[4][3] ),
    .A2(_03521_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09328_ (.A1(_03231_),
    .A2(_03523_),
    .B(_03527_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09329_ (.A1(_03037_),
    .A2(_03519_),
    .B1(_03531_),
    .B2(_03532_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09330_ (.I(_02632_),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09331_ (.A1(\as2650.stack[4][4] ),
    .A2(_03521_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09332_ (.A1(_02456_),
    .A2(_03523_),
    .B(_03527_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09333_ (.A1(_03040_),
    .A2(_03533_),
    .B1(_03534_),
    .B2(_03535_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09334_ (.A1(\as2650.stack[4][5] ),
    .A2(_03526_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09335_ (.A1(_02989_),
    .A2(_02634_),
    .B(_03518_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09336_ (.A1(_03044_),
    .A2(_03533_),
    .B1(_03536_),
    .B2(_03537_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09337_ (.A1(\as2650.stack[4][6] ),
    .A2(_03526_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09338_ (.A1(_03239_),
    .A2(_02634_),
    .B(_03518_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09339_ (.A1(_03047_),
    .A2(_03533_),
    .B1(_03538_),
    .B2(_03539_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09340_ (.A1(\as2650.stack[4][7] ),
    .A2(_03526_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09341_ (.A1(_02129_),
    .A2(_02634_),
    .B(_03518_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09342_ (.A1(_03050_),
    .A2(_03533_),
    .B1(_03540_),
    .B2(_03541_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09343_ (.I(_01030_),
    .Z(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09344_ (.I(_02650_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09345_ (.I(_03543_),
    .Z(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09346_ (.A1(_02143_),
    .A2(_02437_),
    .A3(_02147_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09347_ (.I(_03545_),
    .Z(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09348_ (.A1(\as2650.stack[3][0] ),
    .A2(_03546_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09349_ (.I(_02644_),
    .Z(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09350_ (.A1(_02045_),
    .A2(_03548_),
    .B(_02659_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09351_ (.A1(_03542_),
    .A2(_03544_),
    .B1(_03547_),
    .B2(_03549_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09352_ (.I(_02049_),
    .Z(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09353_ (.A1(_02284_),
    .A2(_02658_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09354_ (.I(_03545_),
    .Z(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09355_ (.I(_02651_),
    .Z(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09356_ (.A1(\as2650.stack[3][1] ),
    .A2(_03552_),
    .B(_03553_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09357_ (.A1(_03550_),
    .A2(_03544_),
    .B1(_03551_),
    .B2(_03554_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09358_ (.I(_02066_),
    .Z(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09359_ (.A1(\as2650.stack[3][2] ),
    .A2(_03546_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09360_ (.A1(_02074_),
    .A2(_03548_),
    .B(_03553_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09361_ (.A1(_03555_),
    .A2(_03544_),
    .B1(_03556_),
    .B2(_03557_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09362_ (.I(_02076_),
    .Z(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09363_ (.A1(\as2650.stack[3][3] ),
    .A2(_03546_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09364_ (.A1(_03231_),
    .A2(_03548_),
    .B(_03553_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09365_ (.A1(_03558_),
    .A2(_03544_),
    .B1(_03559_),
    .B2(_03560_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09366_ (.I(_02090_),
    .Z(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09367_ (.I(_02651_),
    .Z(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09368_ (.A1(\as2650.stack[3][4] ),
    .A2(_03546_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09369_ (.A1(_02456_),
    .A2(_03548_),
    .B(_03553_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09370_ (.A1(_03561_),
    .A2(_03562_),
    .B1(_03563_),
    .B2(_03564_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09371_ (.I(_02100_),
    .Z(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09372_ (.A1(\as2650.stack[3][5] ),
    .A2(_03552_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09373_ (.A1(_02110_),
    .A2(_02653_),
    .B(_03543_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09374_ (.A1(_03565_),
    .A2(_03562_),
    .B1(_03566_),
    .B2(_03567_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09375_ (.I(_02112_),
    .Z(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09376_ (.A1(\as2650.stack[3][6] ),
    .A2(_03552_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09377_ (.A1(_03239_),
    .A2(_02653_),
    .B(_03543_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09378_ (.A1(_03568_),
    .A2(_03562_),
    .B1(_03569_),
    .B2(_03570_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09379_ (.I(_02121_),
    .Z(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09380_ (.A1(\as2650.stack[3][7] ),
    .A2(_03552_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09381_ (.A1(_02129_),
    .A2(_02653_),
    .B(_03543_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09382_ (.A1(_03571_),
    .A2(_03562_),
    .B1(_03572_),
    .B2(_03573_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09383_ (.I(_02510_),
    .Z(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09384_ (.I(_03574_),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09385_ (.A1(_02272_),
    .A2(_03024_),
    .A3(_03218_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09386_ (.I(_03576_),
    .Z(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09387_ (.A1(\as2650.stack[6][0] ),
    .A2(_03577_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09388_ (.I(_02506_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09389_ (.A1(_02045_),
    .A2(_03579_),
    .B(_02523_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09390_ (.A1(_03542_),
    .A2(_03575_),
    .B1(_03578_),
    .B2(_03580_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09391_ (.A1(\as2650.stack[6][1] ),
    .A2(_03577_),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09392_ (.I(_02511_),
    .Z(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09393_ (.A1(_02364_),
    .A2(_03579_),
    .B(_03582_),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09394_ (.A1(_03550_),
    .A2(_03575_),
    .B1(_03581_),
    .B2(_03583_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09395_ (.A1(_02167_),
    .A2(_02522_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09396_ (.I(_03576_),
    .Z(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09397_ (.A1(\as2650.stack[6][2] ),
    .A2(_03585_),
    .B(_03582_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09398_ (.A1(_03555_),
    .A2(_03575_),
    .B1(_03584_),
    .B2(_03586_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09399_ (.A1(\as2650.stack[6][3] ),
    .A2(_03577_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09400_ (.A1(_02087_),
    .A2(_02514_),
    .B(_03582_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09401_ (.A1(_03558_),
    .A2(_03575_),
    .B1(_03587_),
    .B2(_03588_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09402_ (.I(_02511_),
    .Z(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09403_ (.A1(_03509_),
    .A2(_03579_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09404_ (.A1(\as2650.stack[6][4] ),
    .A2(_03585_),
    .B(_03582_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09405_ (.A1(_03561_),
    .A2(_03589_),
    .B1(_03590_),
    .B2(_03591_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09406_ (.A1(_02177_),
    .A2(_03579_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09407_ (.A1(\as2650.stack[6][5] ),
    .A2(_03585_),
    .B(_03574_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09408_ (.A1(_03565_),
    .A2(_03589_),
    .B1(_03592_),
    .B2(_03593_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09409_ (.A1(\as2650.stack[6][6] ),
    .A2(_03577_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09410_ (.A1(_02119_),
    .A2(_02514_),
    .B(_03574_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09411_ (.A1(_03568_),
    .A2(_03589_),
    .B1(_03594_),
    .B2(_03595_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09412_ (.A1(\as2650.stack[6][7] ),
    .A2(_03585_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09413_ (.A1(_02129_),
    .A2(_02514_),
    .B(_03574_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09414_ (.A1(_03571_),
    .A2(_03589_),
    .B1(_03596_),
    .B2(_03597_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09415_ (.A1(_02730_),
    .A2(_02580_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09416_ (.A1(_00677_),
    .A2(_00921_),
    .A3(_00883_),
    .A4(_00768_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09417_ (.A1(_03598_),
    .A2(_03599_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09418_ (.I(_03600_),
    .Z(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09419_ (.I0(\as2650.ivec[0] ),
    .I1(_01102_),
    .S(_03601_),
    .Z(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09420_ (.I(_03602_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09421_ (.I0(\as2650.ivec[1] ),
    .I1(_03261_),
    .S(_03601_),
    .Z(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09422_ (.I(_03603_),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09423_ (.I(_03600_),
    .Z(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09424_ (.I0(\as2650.ivec[2] ),
    .I1(_03267_),
    .S(_03604_),
    .Z(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09425_ (.I(_03605_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09426_ (.I0(\as2650.ivec[3] ),
    .I1(_03273_),
    .S(_03604_),
    .Z(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09427_ (.I(_03606_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09428_ (.I0(\as2650.ivec[4] ),
    .I1(_03279_),
    .S(_03604_),
    .Z(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09429_ (.I(_03607_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09430_ (.I0(\as2650.ivec[5] ),
    .I1(_03285_),
    .S(_03604_),
    .Z(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09431_ (.I(_03608_),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09432_ (.I(_01975_),
    .Z(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09433_ (.I0(\as2650.ivec[6] ),
    .I1(_03609_),
    .S(_03600_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09434_ (.I(_03610_),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09435_ (.A1(\as2650.ivec[7] ),
    .A2(_03601_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09436_ (.A1(_01980_),
    .A2(_03601_),
    .B(_03611_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09437_ (.I(_02533_),
    .Z(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09438_ (.I(_03612_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09439_ (.A1(_02003_),
    .A2(_03024_),
    .A3(_03218_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09440_ (.I(_03614_),
    .Z(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09441_ (.A1(\as2650.stack[5][0] ),
    .A2(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09442_ (.I(_02529_),
    .Z(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09443_ (.A1(_02045_),
    .A2(_03617_),
    .B(_02542_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09444_ (.A1(_03542_),
    .A2(_03613_),
    .B1(_03616_),
    .B2(_03618_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09445_ (.A1(_02284_),
    .A2(_02541_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09446_ (.I(_03614_),
    .Z(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09447_ (.I(_02534_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09448_ (.A1(\as2650.stack[5][1] ),
    .A2(_03620_),
    .B(_03621_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09449_ (.A1(_03550_),
    .A2(_03613_),
    .B1(_03619_),
    .B2(_03622_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09450_ (.A1(\as2650.stack[5][2] ),
    .A2(_03615_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09451_ (.A1(_02074_),
    .A2(_03617_),
    .B(_03621_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09452_ (.A1(_03555_),
    .A2(_03613_),
    .B1(_03623_),
    .B2(_03624_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09453_ (.A1(\as2650.stack[5][3] ),
    .A2(_03615_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09454_ (.A1(_02087_),
    .A2(_02536_),
    .B(_03621_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09455_ (.A1(_03558_),
    .A2(_03613_),
    .B1(_03625_),
    .B2(_03626_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09456_ (.I(_02534_),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09457_ (.A1(_03509_),
    .A2(_03617_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09458_ (.A1(\as2650.stack[5][4] ),
    .A2(_03620_),
    .B(_03621_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09459_ (.A1(_03561_),
    .A2(_03627_),
    .B1(_03628_),
    .B2(_03629_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09460_ (.A1(\as2650.stack[5][5] ),
    .A2(_03615_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09461_ (.A1(_02110_),
    .A2(_02536_),
    .B(_03612_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09462_ (.A1(_03565_),
    .A2(_03627_),
    .B1(_03630_),
    .B2(_03631_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09463_ (.A1(\as2650.stack[5][6] ),
    .A2(_03620_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09464_ (.A1(_02119_),
    .A2(_02536_),
    .B(_03612_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09465_ (.A1(_03568_),
    .A2(_03627_),
    .B1(_03632_),
    .B2(_03633_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09466_ (.A1(_02184_),
    .A2(_03617_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09467_ (.A1(\as2650.stack[5][7] ),
    .A2(_03620_),
    .B(_03612_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09468_ (.A1(_03571_),
    .A2(_03627_),
    .B1(_03634_),
    .B2(_03635_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09469_ (.I(net26),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09470_ (.A1(_00899_),
    .A2(_00758_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09471_ (.I(_00616_),
    .Z(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09472_ (.I(_03638_),
    .Z(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09473_ (.A1(_00622_),
    .A2(_00687_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09474_ (.I(_02823_),
    .Z(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09475_ (.I(_03641_),
    .Z(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09476_ (.A1(_03639_),
    .A2(_03640_),
    .B(_03642_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09477_ (.A1(_00928_),
    .A2(_00772_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09478_ (.A1(_00564_),
    .A2(_03644_),
    .Z(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09479_ (.I(_00541_),
    .Z(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09480_ (.A1(_03646_),
    .A2(_02759_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09481_ (.A1(_02806_),
    .A2(_03647_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09482_ (.I(_03648_),
    .Z(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09483_ (.I(_00973_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09484_ (.A1(_02732_),
    .A2(_03650_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09485_ (.A1(_00465_),
    .A2(_03645_),
    .B1(_03649_),
    .B2(_03651_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09486_ (.A1(_00502_),
    .A2(_00504_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09487_ (.A1(_00879_),
    .A2(_02348_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09488_ (.A1(_00773_),
    .A2(_00785_),
    .A3(_03654_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09489_ (.A1(_02566_),
    .A2(_01712_),
    .B(_02761_),
    .C(_03655_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09490_ (.I(_00504_),
    .Z(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09491_ (.A1(_03657_),
    .A2(_02546_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09492_ (.A1(_02568_),
    .A2(_03653_),
    .A3(_03656_),
    .A4(_03658_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09493_ (.A1(_03637_),
    .A2(_03643_),
    .B(_03652_),
    .C(_03659_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09494_ (.I(_02807_),
    .Z(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09495_ (.I(_03661_),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09496_ (.A1(_02809_),
    .A2(_00694_),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09497_ (.A1(_03662_),
    .A2(_00623_),
    .B(_03660_),
    .C(_03663_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09498_ (.A1(_03636_),
    .A2(_03660_),
    .B(_03664_),
    .C(_00697_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09499_ (.I(_00929_),
    .Z(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09500_ (.A1(_03665_),
    .A2(_03638_),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09501_ (.I(_03666_),
    .Z(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09502_ (.A1(_00825_),
    .A2(_02352_),
    .B(_00648_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09503_ (.A1(_00901_),
    .A2(_02555_),
    .A3(_03667_),
    .A4(_03668_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09504_ (.A1(net24),
    .A2(_03669_),
    .B(_02894_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09505_ (.A1(_01091_),
    .A2(_03669_),
    .B(_03670_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09506_ (.I(net25),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09507_ (.A1(_00483_),
    .A2(_02554_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09508_ (.I(_02581_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09509_ (.A1(_00572_),
    .A2(_02553_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09510_ (.A1(_00622_),
    .A2(_00911_),
    .B(_03640_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09511_ (.A1(_00496_),
    .A2(_02548_),
    .A3(_03675_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09512_ (.A1(_03674_),
    .A2(_03676_),
    .Z(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09513_ (.A1(_02823_),
    .A2(_02568_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09514_ (.I(_03653_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09515_ (.A1(_00865_),
    .A2(_00787_),
    .A3(_03678_),
    .A4(_03679_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09516_ (.A1(_00648_),
    .A2(_02593_),
    .B(_03680_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09517_ (.A1(_02726_),
    .A2(_03673_),
    .B(_03677_),
    .C(_03681_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09518_ (.I0(_03671_),
    .I1(_03672_),
    .S(_03682_),
    .Z(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09519_ (.A1(_02625_),
    .A2(_03683_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09520_ (.A1(_00442_),
    .A2(_00782_),
    .A3(_02737_),
    .A4(_03672_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09521_ (.A1(_02552_),
    .A2(_00547_),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09522_ (.A1(_01005_),
    .A2(_00905_),
    .A3(_00986_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09523_ (.A1(_00985_),
    .A2(_03685_),
    .A3(_03686_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09524_ (.A1(_00616_),
    .A2(_02593_),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09525_ (.A1(_00772_),
    .A2(_00784_),
    .A3(_01712_),
    .A4(_02580_),
    .Z(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09526_ (.A1(_03688_),
    .A2(_03689_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09527_ (.A1(_00577_),
    .A2(_00579_),
    .A3(_00581_),
    .B(_00567_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09528_ (.I(_02017_),
    .Z(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09529_ (.A1(_02599_),
    .A2(_03691_),
    .B(_02549_),
    .C(_03692_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09530_ (.A1(_00878_),
    .A2(_00490_),
    .A3(_00669_),
    .A4(_02550_),
    .Z(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09531_ (.A1(_00832_),
    .A2(_02567_),
    .A3(_02738_),
    .B1(_03694_),
    .B2(_00778_),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09532_ (.A1(_05697_),
    .A2(_00840_),
    .A3(_00870_),
    .A4(_02555_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09533_ (.A1(_02585_),
    .A2(_02578_),
    .A3(_03695_),
    .A4(_03696_),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09534_ (.A1(_03687_),
    .A2(_03690_),
    .A3(_03693_),
    .A4(_03697_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09535_ (.A1(_00852_),
    .A2(_02588_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09536_ (.A1(_02563_),
    .A2(_03699_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09537_ (.A1(_02594_),
    .A2(_02602_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09538_ (.A1(_00467_),
    .A2(_02016_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09539_ (.A1(_00901_),
    .A2(_02004_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09540_ (.A1(_03702_),
    .A2(_03703_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09541_ (.A1(_00891_),
    .A2(_02005_),
    .A3(_02572_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09542_ (.A1(_00735_),
    .A2(_00729_),
    .B(_03704_),
    .C(_03705_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09543_ (.A1(_00747_),
    .A2(_00546_),
    .A3(_03645_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09544_ (.A1(_05703_),
    .A2(_00458_),
    .A3(_00949_),
    .A4(_03672_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09545_ (.A1(_02556_),
    .A2(_03708_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09546_ (.A1(_03707_),
    .A2(_03709_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09547_ (.I(_03710_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09548_ (.A1(_00703_),
    .A2(_01712_),
    .A3(_02580_),
    .Z(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09549_ (.A1(_00911_),
    .A2(_00574_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09550_ (.A1(_02552_),
    .A2(_03713_),
    .A3(_00607_),
    .A4(_00956_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09551_ (.A1(_03711_),
    .A2(_03712_),
    .A3(_03714_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09552_ (.A1(_02581_),
    .A2(_02584_),
    .B(_02561_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09553_ (.A1(_03701_),
    .A2(_03706_),
    .A3(_03715_),
    .A4(_03716_),
    .Z(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09554_ (.A1(_03684_),
    .A2(_03698_),
    .A3(_03700_),
    .A4(_03717_),
    .Z(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09555_ (.I(_03718_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09556_ (.I(_03719_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09557_ (.I(_03720_),
    .Z(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09558_ (.I(_02037_),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09559_ (.I(_03722_),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09560_ (.A1(_00748_),
    .A2(_02866_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09561_ (.I(_03724_),
    .Z(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09562_ (.I(_02039_),
    .Z(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09563_ (.A1(_00804_),
    .A2(_02865_),
    .A3(_00816_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09564_ (.I(_03727_),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09565_ (.A1(net90),
    .A2(net8),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09566_ (.A1(_02037_),
    .A2(_01041_),
    .Z(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09567_ (.A1(_03729_),
    .A2(_03730_),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09568_ (.I(net93),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09569_ (.I(_00793_),
    .Z(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09570_ (.I(_03733_),
    .Z(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09571_ (.A1(_03732_),
    .A2(_03734_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09572_ (.A1(_00795_),
    .A2(_03731_),
    .B(_03735_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09573_ (.I(_00672_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09574_ (.A1(_03723_),
    .A2(_05672_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09575_ (.I(_01042_),
    .Z(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09576_ (.I(_03739_),
    .Z(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09577_ (.A1(_00638_),
    .A2(_00893_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09578_ (.I(_03741_),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09579_ (.I(_00681_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09580_ (.I(_03743_),
    .Z(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09581_ (.I(_01130_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09582_ (.I(_03745_),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09583_ (.A1(_03732_),
    .A2(_03744_),
    .B(_03746_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09584_ (.A1(_03740_),
    .A2(_00683_),
    .B1(_03742_),
    .B2(_03732_),
    .C(_03747_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09585_ (.I(_02865_),
    .Z(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09586_ (.I(_00778_),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09587_ (.A1(_03750_),
    .A2(_02747_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09588_ (.I(_03751_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09589_ (.A1(_03749_),
    .A2(_03752_),
    .B(_03723_),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09590_ (.A1(_03737_),
    .A2(_03738_),
    .B1(_03748_),
    .B2(_03753_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09591_ (.I(_00799_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09592_ (.A1(_03728_),
    .A2(_03736_),
    .B(_03754_),
    .C(_03755_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09593_ (.A1(_02745_),
    .A2(_00748_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09594_ (.A1(_03726_),
    .A2(_00801_),
    .B(_03756_),
    .C(_03757_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09595_ (.I(_00538_),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09596_ (.I(_00722_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09597_ (.I(_03760_),
    .Z(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09598_ (.I(_01128_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09599_ (.I(_03762_),
    .Z(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09600_ (.A1(_03740_),
    .A2(_03763_),
    .A3(_01018_),
    .Z(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09601_ (.A1(_03763_),
    .A2(_01019_),
    .B(_03740_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09602_ (.I(_00991_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09603_ (.A1(_03766_),
    .A2(_03092_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09604_ (.A1(_02844_),
    .A2(_03767_),
    .Z(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09605_ (.I(_01005_),
    .Z(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09606_ (.A1(_03761_),
    .A2(_03764_),
    .A3(_03765_),
    .B1(_03768_),
    .B2(_03769_),
    .ZN(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09607_ (.A1(_00538_),
    .A2(_00723_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09608_ (.I(_03771_),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09609_ (.I(net93),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09610_ (.I(_00551_),
    .Z(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09611_ (.A1(_03759_),
    .A2(_03770_),
    .B1(_03772_),
    .B2(_03773_),
    .C(_03774_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09612_ (.I(_00632_),
    .Z(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09613_ (.I(_03776_),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09614_ (.A1(_03777_),
    .A2(_03731_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09615_ (.I(_00730_),
    .Z(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09616_ (.I(_03779_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09617_ (.I(_03654_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09618_ (.I(_03781_),
    .Z(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09619_ (.A1(_03775_),
    .A2(_03778_),
    .B(_03780_),
    .C(_03782_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09620_ (.A1(_03723_),
    .A2(_03725_),
    .B(_03758_),
    .C(_03783_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09621_ (.A1(_03732_),
    .A2(_03720_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09622_ (.I(_00696_),
    .Z(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09623_ (.A1(_03721_),
    .A2(_03784_),
    .B(_03785_),
    .C(_03786_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09624_ (.I(_02055_),
    .Z(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09625_ (.I(_03724_),
    .Z(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09626_ (.I(_00552_),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09627_ (.I(net9),
    .Z(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09628_ (.A1(_02054_),
    .A2(_03790_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09629_ (.A1(_03730_),
    .A2(_03791_),
    .Z(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09630_ (.I(_00538_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09631_ (.I(_03760_),
    .Z(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09632_ (.I(net9),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09633_ (.I(_03795_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09634_ (.I(_03796_),
    .Z(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09635_ (.A1(_01041_),
    .A2(_01018_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09636_ (.A1(_03796_),
    .A2(_01118_),
    .A3(_01158_),
    .Z(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09637_ (.A1(_03798_),
    .A2(_03799_),
    .Z(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09638_ (.A1(_03762_),
    .A2(_03800_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09639_ (.A1(_03797_),
    .A2(_03763_),
    .B(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09640_ (.I(_03766_),
    .Z(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09641_ (.A1(_01041_),
    .A2(_03092_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09642_ (.A1(_03796_),
    .A2(_01118_),
    .A3(_01124_),
    .Z(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09643_ (.A1(_03804_),
    .A2(_03805_),
    .B(_01002_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09644_ (.A1(_03804_),
    .A2(_03805_),
    .B(_03806_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09645_ (.A1(_03797_),
    .A2(_03803_),
    .B(_03807_),
    .C(_00534_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09646_ (.A1(_03794_),
    .A2(_03802_),
    .B(_03808_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09647_ (.A1(net31),
    .A2(_03773_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09648_ (.I(_03771_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09649_ (.A1(_03793_),
    .A2(_03809_),
    .B1(_03810_),
    .B2(_03811_),
    .C(_00552_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09650_ (.I(_02889_),
    .Z(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09651_ (.A1(_03789_),
    .A2(_03792_),
    .B(_03812_),
    .C(_03813_),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09652_ (.I(_03657_),
    .Z(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09653_ (.I(_02608_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09654_ (.A1(_00805_),
    .A2(_00816_),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09655_ (.A1(_03816_),
    .A2(_03817_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09656_ (.I(net31),
    .Z(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09657_ (.I(_02952_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09658_ (.A1(_03729_),
    .A2(_03791_),
    .Z(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09659_ (.A1(_00629_),
    .A2(_03821_),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09660_ (.A1(_03819_),
    .A2(_03820_),
    .B(_03822_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09661_ (.I(_03743_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09662_ (.A1(_03824_),
    .A2(_03810_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09663_ (.A1(_02846_),
    .A2(_00683_),
    .B1(_03742_),
    .B2(_03819_),
    .C(_03825_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09664_ (.A1(_02582_),
    .A2(_00815_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09665_ (.A1(_02332_),
    .A2(_03752_),
    .B(_03787_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09666_ (.A1(_03818_),
    .A2(_03823_),
    .B1(_03826_),
    .B2(_03827_),
    .C(_03828_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09667_ (.I(_00451_),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09668_ (.A1(_03787_),
    .A2(_03815_),
    .B1(_03829_),
    .B2(_03830_),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09669_ (.I(_03779_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09670_ (.A1(_03814_),
    .A2(_03831_),
    .B(_03832_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09671_ (.A1(_03787_),
    .A2(_03788_),
    .B(_03833_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09672_ (.A1(_03819_),
    .A2(_03720_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09673_ (.A1(_03721_),
    .A2(_03834_),
    .B(_03835_),
    .C(_03786_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09674_ (.I(net32),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09675_ (.I(_03719_),
    .Z(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09676_ (.A1(net89),
    .A2(net10),
    .Z(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09677_ (.A1(_02055_),
    .A2(_01141_),
    .Z(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09678_ (.A1(_03730_),
    .A2(_03791_),
    .B(_03839_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09679_ (.A1(_03838_),
    .A2(_03840_),
    .Z(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _09680_ (.A1(_03796_),
    .A2(_01125_),
    .A3(_01126_),
    .B1(_03804_),
    .B2(_03805_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09681_ (.A1(_01254_),
    .A2(_01258_),
    .A3(_01260_),
    .B(_01273_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09682_ (.A1(_02849_),
    .A2(_01261_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09683_ (.A1(_03843_),
    .A2(_03844_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09684_ (.A1(_03842_),
    .A2(_03845_),
    .B(_01002_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09685_ (.A1(_03842_),
    .A2(_03845_),
    .B(_03846_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09686_ (.A1(_02850_),
    .A2(_03803_),
    .B(_03847_),
    .C(_00533_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09687_ (.I(_00980_),
    .Z(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09688_ (.I(_03849_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _09689_ (.A1(_03797_),
    .A2(_01159_),
    .A3(_01160_),
    .B1(_03798_),
    .B2(_03799_),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09690_ (.A1(_02848_),
    .A2(_01286_),
    .A3(_03851_),
    .Z(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09691_ (.A1(_01274_),
    .A2(_03849_),
    .B(_03760_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09692_ (.A1(_03850_),
    .A2(_03852_),
    .B(_03853_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09693_ (.A1(_03848_),
    .A2(_03854_),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09694_ (.A1(_03819_),
    .A2(net93),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09695_ (.A1(_03836_),
    .A2(_03856_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09696_ (.A1(_03793_),
    .A2(_03855_),
    .B1(_03857_),
    .B2(_03771_),
    .C(_00551_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09697_ (.I(_02889_),
    .Z(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09698_ (.A1(_03774_),
    .A2(_03841_),
    .B(_03858_),
    .C(_03859_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09699_ (.A1(_02070_),
    .A2(_01271_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09700_ (.A1(_02054_),
    .A2(_03790_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09701_ (.A1(_02054_),
    .A2(_03790_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09702_ (.A1(_03729_),
    .A2(_03862_),
    .B(_03863_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09703_ (.A1(_03861_),
    .A2(_03864_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09704_ (.I(_02932_),
    .Z(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09705_ (.I(_03866_),
    .Z(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09706_ (.A1(_03836_),
    .A2(_03867_),
    .B(_00679_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09707_ (.A1(_00630_),
    .A2(_03865_),
    .B(_03868_),
    .C(_03728_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09708_ (.I(_00638_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09709_ (.A1(_03870_),
    .A2(_03743_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09710_ (.I(_03871_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09711_ (.I(_03744_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _09712_ (.A1(_02851_),
    .A2(_03872_),
    .B1(_03857_),
    .B2(_03873_),
    .C1(_00818_),
    .C2(_03836_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09713_ (.A1(_00523_),
    .A2(_03827_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09714_ (.I(net89),
    .Z(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09715_ (.I(_02607_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09716_ (.A1(_03665_),
    .A2(_03877_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09717_ (.A1(_03752_),
    .A2(_03878_),
    .ZN(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09718_ (.A1(_03876_),
    .A2(_02808_),
    .A3(_03879_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09719_ (.A1(_03874_),
    .A2(_03875_),
    .B(_03880_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09720_ (.A1(_03860_),
    .A2(_03869_),
    .A3(_03881_),
    .B(_00731_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09721_ (.I(_03718_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09722_ (.A1(_02071_),
    .A2(_03725_),
    .B(_03882_),
    .C(_03883_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09723_ (.A1(_03836_),
    .A2(_03837_),
    .B(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09724_ (.A1(_00728_),
    .A2(_03885_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09725_ (.I(net33),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09726_ (.I(_01002_),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09727_ (.I(_03887_),
    .Z(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09728_ (.A1(_01273_),
    .A2(_01254_),
    .A3(_01258_),
    .A4(_01260_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09729_ (.A1(_03842_),
    .A2(_03843_),
    .B(_03889_),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09730_ (.A1(_02854_),
    .A2(_01303_),
    .A3(_03890_),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09731_ (.A1(_03887_),
    .A2(_03891_),
    .B(_00533_),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09732_ (.A1(_02856_),
    .A2(_03888_),
    .B(_03892_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09733_ (.I(_03762_),
    .Z(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09734_ (.A1(_01281_),
    .A2(_01283_),
    .A3(_01285_),
    .B(_01273_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09735_ (.A1(_01272_),
    .A2(_01281_),
    .A3(_01283_),
    .A4(_01285_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09736_ (.A1(_03851_),
    .A2(_03895_),
    .B(_03896_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09737_ (.A1(_02854_),
    .A2(_01322_),
    .A3(_03897_),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09738_ (.A1(_03150_),
    .A2(_03762_),
    .B(_00641_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09739_ (.A1(_03894_),
    .A2(_03898_),
    .B(_03899_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09740_ (.A1(_03893_),
    .A2(_03900_),
    .B(_03793_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09741_ (.A1(net32),
    .A2(net31),
    .A3(net93),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09742_ (.A1(_03886_),
    .A2(_03902_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09743_ (.A1(_03811_),
    .A2(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09744_ (.A1(_00633_),
    .A2(_03901_),
    .A3(_03904_),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09745_ (.A1(_02080_),
    .A2(net11),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09746_ (.A1(_02081_),
    .A2(_01310_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09747_ (.A1(_03906_),
    .A2(_03907_),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09748_ (.A1(_03876_),
    .A2(net10),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09749_ (.A1(_03861_),
    .A2(_03840_),
    .B(_03909_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09750_ (.A1(_03908_),
    .A2(_03910_),
    .B(_03776_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09751_ (.A1(_03908_),
    .A2(_03910_),
    .B(_03911_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09752_ (.A1(_00731_),
    .A2(_03782_),
    .A3(_03905_),
    .A4(_03912_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09753_ (.I(_02080_),
    .Z(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09754_ (.A1(_00881_),
    .A2(_00730_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09755_ (.I(_03915_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09756_ (.I(_03817_),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09757_ (.I(_03909_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09758_ (.A1(_03838_),
    .A2(_03864_),
    .B(_03918_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09759_ (.A1(_03908_),
    .A2(_03919_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09760_ (.I(_01697_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09761_ (.A1(_03886_),
    .A2(_03921_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09762_ (.A1(_03734_),
    .A2(_03920_),
    .B(_03922_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09763_ (.A1(_02855_),
    .A2(_00683_),
    .B1(_03742_),
    .B2(_03886_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09764_ (.I(_00704_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09765_ (.A1(_00689_),
    .A2(_03903_),
    .B(_03924_),
    .C(_03925_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09766_ (.A1(_03917_),
    .A2(_03923_),
    .B(_03926_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09767_ (.A1(_02082_),
    .A2(_03879_),
    .B1(_03927_),
    .B2(_03878_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09768_ (.A1(_03914_),
    .A2(_03725_),
    .B1(_03916_),
    .B2(_03928_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09769_ (.A1(_03913_),
    .A2(_03929_),
    .B(_03883_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09770_ (.A1(_03886_),
    .A2(_03837_),
    .B(_03930_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09771_ (.A1(_00728_),
    .A2(_03931_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09772_ (.A1(_02093_),
    .A2(net12),
    .Z(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09773_ (.I(_03932_),
    .Z(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09774_ (.A1(_03907_),
    .A2(_03910_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09775_ (.A1(_03906_),
    .A2(_03934_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09776_ (.A1(_03933_),
    .A2(_03935_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09777_ (.A1(_02853_),
    .A2(_01302_),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09778_ (.A1(_02852_),
    .A2(_01302_),
    .B1(_03842_),
    .B2(_03843_),
    .C(_03889_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09779_ (.A1(_03937_),
    .A2(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09780_ (.A1(_02858_),
    .A2(_01429_),
    .A3(_03939_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09781_ (.A1(_03888_),
    .A2(_03940_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09782_ (.A1(_02859_),
    .A2(_03803_),
    .B(_00534_),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09783_ (.A1(_02853_),
    .A2(_03147_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09784_ (.A1(_02852_),
    .A2(_03147_),
    .B1(_03851_),
    .B2(_03895_),
    .C(_03896_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09785_ (.A1(_03943_),
    .A2(_03944_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09786_ (.A1(_03165_),
    .A2(_01445_),
    .A3(_03945_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09787_ (.A1(_03763_),
    .A2(_03946_),
    .ZN(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09788_ (.I(_00641_),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09789_ (.A1(_02859_),
    .A2(_03894_),
    .B(_03947_),
    .C(_03948_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09790_ (.A1(_03941_),
    .A2(_03942_),
    .B(_03949_),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09791_ (.I(net34),
    .Z(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09792_ (.I(net33),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09793_ (.A1(_03952_),
    .A2(_03902_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09794_ (.A1(_03951_),
    .A2(_03953_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09795_ (.A1(_03759_),
    .A2(_03950_),
    .B1(_03954_),
    .B2(_03772_),
    .C(_03789_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09796_ (.A1(_00717_),
    .A2(_03936_),
    .B(_03955_),
    .C(_02890_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09797_ (.I(net60),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09798_ (.I(_03957_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09799_ (.I(_03879_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09800_ (.I(_00688_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _09801_ (.A1(_02859_),
    .A2(_03872_),
    .B1(_03954_),
    .B2(_03960_),
    .C1(_00818_),
    .C2(_03951_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09802_ (.A1(_03838_),
    .A2(_03864_),
    .B(_03907_),
    .C(_03918_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09803_ (.A1(_03906_),
    .A2(_03962_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09804_ (.A1(_03933_),
    .A2(_03963_),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09805_ (.A1(_00629_),
    .A2(_03964_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09806_ (.A1(_03951_),
    .A2(_03867_),
    .B(_03965_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09807_ (.A1(_00816_),
    .A2(_03961_),
    .B1(_03966_),
    .B2(_03917_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09808_ (.I(_03878_),
    .Z(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09809_ (.A1(_03958_),
    .A2(_03959_),
    .B1(_03967_),
    .B2(_03968_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09810_ (.A1(_02094_),
    .A2(_03725_),
    .B1(_03916_),
    .B2(_03969_),
    .C(_03883_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09811_ (.A1(_00822_),
    .A2(_03956_),
    .B(_03970_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09812_ (.I(_02893_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09813_ (.A1(_03951_),
    .A2(_03837_),
    .B(_03972_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09814_ (.A1(_03971_),
    .A2(_03973_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09815_ (.I(_00727_),
    .Z(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09816_ (.I(net35),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09817_ (.I(_03719_),
    .Z(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09818_ (.I(_00748_),
    .Z(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09819_ (.I(_01434_),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09820_ (.A1(_03978_),
    .A2(_01428_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09821_ (.A1(_03978_),
    .A2(_01428_),
    .ZN(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09822_ (.A1(_03937_),
    .A2(_03979_),
    .A3(_03938_),
    .B(_03980_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09823_ (.A1(_01466_),
    .A2(_01458_),
    .A3(_03981_),
    .Z(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09824_ (.A1(_03803_),
    .A2(_03982_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09825_ (.A1(_02613_),
    .A2(_03887_),
    .B(_01005_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09826_ (.A1(_03978_),
    .A2(_01444_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09827_ (.A1(_03978_),
    .A2(_01444_),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09828_ (.A1(_03943_),
    .A2(_03985_),
    .A3(_03944_),
    .B(_03986_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09829_ (.A1(_02612_),
    .A2(_01474_),
    .Z(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09830_ (.A1(_03987_),
    .A2(_03988_),
    .B(_03849_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09831_ (.A1(_03987_),
    .A2(_03988_),
    .B(_03989_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09832_ (.I(_03760_),
    .Z(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09833_ (.A1(_02612_),
    .A2(_03850_),
    .B(_03991_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09834_ (.A1(_03983_),
    .A2(_03984_),
    .B1(_03990_),
    .B2(_03992_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09835_ (.A1(_00718_),
    .A2(_03993_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09836_ (.A1(_03793_),
    .A2(_00723_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09837_ (.A1(net34),
    .A2(_03953_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09838_ (.A1(net35),
    .A2(_03996_),
    .Z(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09839_ (.A1(_03995_),
    .A2(_03997_),
    .B(_03776_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09840_ (.A1(_02105_),
    .A2(_01464_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09841_ (.I(_03999_),
    .Z(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09842_ (.A1(_03933_),
    .A2(_03935_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09843_ (.A1(_03958_),
    .A2(_02858_),
    .B(_04001_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09844_ (.A1(_04000_),
    .A2(_04002_),
    .Z(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09845_ (.I(_03776_),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09846_ (.A1(_03994_),
    .A2(_03998_),
    .B1(_04003_),
    .B2(_04004_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09847_ (.A1(_03977_),
    .A2(_02890_),
    .A3(_04005_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09848_ (.I(net61),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09849_ (.A1(_00800_),
    .A2(_02618_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09850_ (.I(_00698_),
    .Z(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09851_ (.A1(_03870_),
    .A2(_02612_),
    .A3(_03743_),
    .Z(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09852_ (.A1(_03975_),
    .A2(_03742_),
    .B1(_03997_),
    .B2(_04009_),
    .C(_04010_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09853_ (.A1(_03975_),
    .A2(_02955_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09854_ (.A1(_03933_),
    .A2(_03963_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09855_ (.A1(_03957_),
    .A2(_01435_),
    .B(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09856_ (.A1(_04000_),
    .A2(_04014_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09857_ (.A1(_00629_),
    .A2(_04015_),
    .B(_03817_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09858_ (.A1(_03925_),
    .A2(_04011_),
    .B1(_04012_),
    .B2(_04016_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09859_ (.A1(_04008_),
    .A2(_04017_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09860_ (.A1(_02107_),
    .A2(_03959_),
    .B(_04018_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09861_ (.A1(_04007_),
    .A2(_03724_),
    .B1(_03916_),
    .B2(_04019_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09862_ (.A1(_04006_),
    .A2(_04020_),
    .B(_03883_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09863_ (.A1(_03975_),
    .A2(_03976_),
    .B(_04021_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09864_ (.A1(_03974_),
    .A2(_04022_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09865_ (.I(_02115_),
    .Z(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09866_ (.I(_00534_),
    .Z(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09867_ (.I(_02826_),
    .Z(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09868_ (.A1(_01609_),
    .A2(_01618_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09869_ (.A1(_01465_),
    .A2(_01457_),
    .Z(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09870_ (.A1(_02611_),
    .A2(_01457_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09871_ (.A1(_03981_),
    .A2(_04027_),
    .B(_04028_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09872_ (.A1(_04026_),
    .A2(_04029_),
    .B(_03766_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09873_ (.A1(_04026_),
    .A2(_04029_),
    .B(_04030_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09874_ (.A1(_04025_),
    .A2(_03888_),
    .B(_04031_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09875_ (.A1(_02861_),
    .A2(_03850_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09876_ (.A1(_01609_),
    .A2(_01596_),
    .Z(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09877_ (.A1(_02611_),
    .A2(_01473_),
    .Z(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09878_ (.A1(_02611_),
    .A2(_01473_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09879_ (.A1(_03987_),
    .A2(_04035_),
    .B(_04036_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09880_ (.A1(_04034_),
    .A2(_04037_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09881_ (.A1(_03894_),
    .A2(_04038_),
    .B(_03794_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09882_ (.A1(_04024_),
    .A2(_04032_),
    .B1(_04033_),
    .B2(_04039_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09883_ (.I(net36),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09884_ (.A1(_03975_),
    .A2(_03996_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09885_ (.A1(_04041_),
    .A2(_04042_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09886_ (.A1(_03811_),
    .A2(_04043_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09887_ (.A1(_00718_),
    .A2(_04040_),
    .B(_04044_),
    .C(_04004_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09888_ (.A1(net62),
    .A2(_01607_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09889_ (.I(_04046_),
    .Z(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09890_ (.A1(net62),
    .A2(_01607_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09891_ (.A1(_04047_),
    .A2(_04048_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09892_ (.A1(_03957_),
    .A2(net12),
    .B1(_01464_),
    .B2(_02105_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09893_ (.A1(_02106_),
    .A2(_02933_),
    .B(_04050_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09894_ (.A1(_04001_),
    .A2(_04000_),
    .B(_04051_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09895_ (.A1(_04049_),
    .A2(_04052_),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09896_ (.A1(_03774_),
    .A2(_04053_),
    .B(_03813_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09897_ (.A1(_04013_),
    .A2(_03999_),
    .B(_04051_),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09898_ (.A1(_04049_),
    .A2(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09899_ (.A1(_04041_),
    .A2(_03820_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09900_ (.A1(_00810_),
    .A2(_04056_),
    .B(_04057_),
    .C(_03917_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09901_ (.A1(_04025_),
    .A2(_03872_),
    .B1(_00817_),
    .B2(_04041_),
    .C(_03925_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09902_ (.A1(_00896_),
    .A2(_04043_),
    .B(_04059_),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09903_ (.A1(_04058_),
    .A2(_04060_),
    .B(_03968_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09904_ (.I(_02745_),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09905_ (.A1(_04023_),
    .A2(_03959_),
    .B(_04062_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09906_ (.A1(_04045_),
    .A2(_04054_),
    .B1(_04061_),
    .B2(_04063_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09907_ (.A1(_04023_),
    .A2(_03788_),
    .B1(_04064_),
    .B2(_03977_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09908_ (.A1(_04041_),
    .A2(_03720_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09909_ (.A1(_03837_),
    .A2(_04065_),
    .B(_04066_),
    .C(_03786_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09910_ (.I(_03719_),
    .Z(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09911_ (.I(_04067_),
    .Z(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09912_ (.I(_03724_),
    .Z(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09913_ (.A1(_01610_),
    .A2(_01619_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09914_ (.A1(_04026_),
    .A2(_04029_),
    .B(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09915_ (.A1(_00808_),
    .A2(_01693_),
    .Z(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09916_ (.A1(_04071_),
    .A2(_04072_),
    .B(_03887_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09917_ (.A1(_04071_),
    .A2(_04072_),
    .B(_04073_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09918_ (.I(_00626_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09919_ (.I(_04075_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09920_ (.I(_04076_),
    .Z(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09921_ (.I(_04077_),
    .Z(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09922_ (.A1(_04078_),
    .A2(_03888_),
    .B(_03769_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09923_ (.A1(_04078_),
    .A2(_03850_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09924_ (.A1(_01592_),
    .A2(_01594_),
    .A3(_01595_),
    .Z(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09925_ (.A1(_01610_),
    .A2(_04081_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09926_ (.A1(_04034_),
    .A2(_04037_),
    .B(_04082_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09927_ (.A1(_04076_),
    .A2(_01696_),
    .A3(_04083_),
    .Z(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09928_ (.A1(_03894_),
    .A2(_04084_),
    .B(_03761_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09929_ (.A1(_04074_),
    .A2(_04079_),
    .B1(_04080_),
    .B2(_04085_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09930_ (.I(net37),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09931_ (.A1(net36),
    .A2(net35),
    .A3(_03996_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09932_ (.A1(_04087_),
    .A2(_04088_),
    .Z(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09933_ (.A1(_03772_),
    .A2(_04089_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09934_ (.A1(_00719_),
    .A2(_04086_),
    .B(_04090_),
    .C(_03777_),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09935_ (.A1(net63),
    .A2(net2),
    .Z(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09936_ (.A1(_04049_),
    .A2(_04052_),
    .B(_04047_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09937_ (.A1(_04092_),
    .A2(_04093_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09938_ (.A1(_00717_),
    .A2(_04094_),
    .B(_02890_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09939_ (.A1(_04049_),
    .A2(_04055_),
    .B(_04047_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09940_ (.A1(_04092_),
    .A2(_04096_),
    .Z(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09941_ (.A1(_04078_),
    .A2(_04097_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09942_ (.I(_03733_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09943_ (.A1(_04087_),
    .A2(_04099_),
    .B(_03728_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09944_ (.I(_03751_),
    .Z(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09945_ (.I(_00688_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09946_ (.I(_00682_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09947_ (.I(_03741_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09948_ (.I(_00957_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09949_ (.A1(_03866_),
    .A2(_04103_),
    .B1(_04104_),
    .B2(_04087_),
    .C(_04105_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09950_ (.A1(_04102_),
    .A2(_04089_),
    .B(_04106_),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09951_ (.A1(_02126_),
    .A2(_04101_),
    .B(_04107_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09952_ (.I(_00672_),
    .Z(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09953_ (.A1(_04098_),
    .A2(_04100_),
    .B1(_04108_),
    .B2(_04109_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09954_ (.A1(_02808_),
    .A2(_04008_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09955_ (.A1(_03830_),
    .A2(_04110_),
    .B1(_04111_),
    .B2(_02126_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09956_ (.A1(_04091_),
    .A2(_04095_),
    .B(_04112_),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09957_ (.A1(_02126_),
    .A2(_04069_),
    .B1(_04113_),
    .B2(_02606_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09958_ (.A1(_04087_),
    .A2(_03976_),
    .B(_02894_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09959_ (.A1(_04068_),
    .A2(_04114_),
    .B(_04115_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09960_ (.I(\as2650.addr_buff[0] ),
    .Z(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09961_ (.A1(_00792_),
    .A2(_01692_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09962_ (.A1(_04026_),
    .A2(_04029_),
    .B(_04117_),
    .C(_04070_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09963_ (.A1(_04075_),
    .A2(_01692_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09964_ (.A1(_00961_),
    .A2(_04119_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09965_ (.A1(_04118_),
    .A2(_04120_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09966_ (.A1(_04116_),
    .A2(_04121_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09967_ (.A1(_04075_),
    .A2(_01695_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09968_ (.A1(_04034_),
    .A2(_04037_),
    .B(_04123_),
    .C(_04082_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09969_ (.A1(_04075_),
    .A2(_01695_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09970_ (.A1(_03849_),
    .A2(_04125_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09971_ (.A1(_04124_),
    .A2(_04126_),
    .ZN(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09972_ (.A1(_04116_),
    .A2(_04127_),
    .Z(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09973_ (.I(_03948_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09974_ (.A1(_04024_),
    .A2(_04122_),
    .B1(_04128_),
    .B2(_04129_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09975_ (.I(net38),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09976_ (.I(net37),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09977_ (.A1(_04132_),
    .A2(_04088_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09978_ (.A1(_04131_),
    .A2(_04133_),
    .Z(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09979_ (.A1(_00719_),
    .A2(_04130_),
    .B1(_04134_),
    .B2(_03995_),
    .C(_03777_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09980_ (.I(_01607_),
    .Z(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09981_ (.A1(net88),
    .A2(_04136_),
    .Z(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09982_ (.A1(_04046_),
    .A2(_04048_),
    .A3(_04092_),
    .Z(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09983_ (.A1(_02125_),
    .A2(_04136_),
    .B1(_04051_),
    .B2(_04138_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09984_ (.A1(_04001_),
    .A2(_04000_),
    .A3(_04138_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09985_ (.A1(_04047_),
    .A2(_04139_),
    .A3(_04140_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09986_ (.A1(_04137_),
    .A2(_04141_),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09987_ (.A1(_04137_),
    .A2(_04141_),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09988_ (.A1(_00633_),
    .A2(_04143_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09989_ (.I(_02889_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09990_ (.A1(_04142_),
    .A2(_04144_),
    .B(_04145_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09991_ (.A1(_04046_),
    .A2(_04139_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09992_ (.A1(_03999_),
    .A2(_04138_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09993_ (.A1(_03932_),
    .A2(_03963_),
    .A3(_04148_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09994_ (.A1(_04147_),
    .A2(_04149_),
    .B(_04137_),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09995_ (.A1(_04137_),
    .A2(_04147_),
    .A3(_04149_),
    .Z(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09996_ (.A1(_04150_),
    .A2(_04151_),
    .Z(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09997_ (.A1(_03734_),
    .A2(_04152_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09998_ (.A1(_04131_),
    .A2(_03867_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09999_ (.A1(_03873_),
    .A2(_04134_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10000_ (.I(\as2650.addr_buff[0] ),
    .Z(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10001_ (.I(_04156_),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10002_ (.A1(_04157_),
    .A2(_03872_),
    .B1(_00818_),
    .B2(_04131_),
    .C(_03925_),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10003_ (.A1(_03917_),
    .A2(_04153_),
    .A3(_04154_),
    .B1(_04155_),
    .B2(_04158_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10004_ (.A1(_02195_),
    .A2(_03959_),
    .B1(_04159_),
    .B2(_03968_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10005_ (.I(_03661_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10006_ (.A1(_04135_),
    .A2(_04146_),
    .B1(_04160_),
    .B2(_04161_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10007_ (.I(_00749_),
    .Z(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10008_ (.A1(_02195_),
    .A2(_04069_),
    .B1(_04162_),
    .B2(_04163_),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10009_ (.I(_02893_),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10010_ (.A1(_04131_),
    .A2(_03976_),
    .B(_04165_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10011_ (.A1(_04068_),
    .A2(_04164_),
    .B(_04166_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10012_ (.I(net87),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10013_ (.A1(_04167_),
    .A2(_04136_),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10014_ (.I(_04168_),
    .Z(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10015_ (.A1(_02193_),
    .A2(_02940_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10016_ (.A1(_04170_),
    .A2(_04142_),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10017_ (.A1(_04169_),
    .A2(_04171_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10018_ (.I(\as2650.addr_buff[1] ),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10019_ (.I(_04173_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10020_ (.I(_04174_),
    .Z(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10021_ (.A1(_04156_),
    .A2(_04124_),
    .A3(_04126_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10022_ (.A1(_04175_),
    .A2(_04176_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10023_ (.A1(_04156_),
    .A2(_04118_),
    .A3(_04120_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10024_ (.A1(_04174_),
    .A2(_04178_),
    .Z(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10025_ (.A1(_03794_),
    .A2(_04177_),
    .B1(_04179_),
    .B2(_03769_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10026_ (.I(net39),
    .Z(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10027_ (.A1(net38),
    .A2(_04133_),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10028_ (.A1(_04181_),
    .A2(_04182_),
    .Z(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10029_ (.A1(_03759_),
    .A2(_04180_),
    .B1(_04183_),
    .B2(_03811_),
    .C(_00552_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10030_ (.A1(_03789_),
    .A2(_04172_),
    .B(_04184_),
    .C(_04145_),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10031_ (.I(_04173_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10032_ (.A1(_04186_),
    .A2(_00682_),
    .B1(_04104_),
    .B2(_04181_),
    .C(_04105_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10033_ (.A1(_03824_),
    .A2(_04183_),
    .B(_04187_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10034_ (.A1(_02205_),
    .A2(_04101_),
    .B(_04188_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10035_ (.A1(_04181_),
    .A2(_04099_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10036_ (.A1(_04170_),
    .A2(_04150_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10037_ (.A1(_04169_),
    .A2(_04191_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10038_ (.A1(_04078_),
    .A2(_04192_),
    .B(_03727_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10039_ (.A1(_04109_),
    .A2(_04189_),
    .B1(_04190_),
    .B2(_04193_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10040_ (.A1(_02205_),
    .A2(_04111_),
    .B1(_04194_),
    .B2(_03830_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10041_ (.A1(_04185_),
    .A2(_04195_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10042_ (.A1(_02205_),
    .A2(_04069_),
    .B1(_04196_),
    .B2(_04163_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10043_ (.A1(_04181_),
    .A2(_03976_),
    .B(_04165_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10044_ (.A1(_04068_),
    .A2(_04197_),
    .B(_04198_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10045_ (.I(\as2650.addr_buff[2] ),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10046_ (.I(_04199_),
    .Z(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10047_ (.A1(_04175_),
    .A2(_04176_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10048_ (.A1(\as2650.addr_buff[0] ),
    .A2(_04173_),
    .A3(\as2650.addr_buff[2] ),
    .Z(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10049_ (.A1(_04124_),
    .A2(_04126_),
    .A3(_04202_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10050_ (.A1(_04200_),
    .A2(_04201_),
    .B(_04203_),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10051_ (.A1(_04175_),
    .A2(_04178_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10052_ (.A1(_04118_),
    .A2(_04120_),
    .A3(_04202_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10053_ (.A1(_04200_),
    .A2(_04205_),
    .B(_04206_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10054_ (.A1(_04129_),
    .A2(_04204_),
    .B1(_04207_),
    .B2(_04024_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10055_ (.I(net40),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10056_ (.A1(net39),
    .A2(net38),
    .A3(_04133_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10057_ (.A1(_04209_),
    .A2(_04210_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10058_ (.A1(_00718_),
    .A2(_04208_),
    .B1(_04211_),
    .B2(_03995_),
    .C(_04004_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10059_ (.A1(_02204_),
    .A2(_01611_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10060_ (.A1(_04170_),
    .A2(_04213_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10061_ (.A1(_04142_),
    .A2(_04169_),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10062_ (.A1(net66),
    .A2(_01608_),
    .Z(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10063_ (.I(_04216_),
    .Z(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10064_ (.A1(_04214_),
    .A2(_04215_),
    .B(_04217_),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10065_ (.A1(_04217_),
    .A2(_04214_),
    .A3(_04215_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10066_ (.A1(_00633_),
    .A2(_04219_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10067_ (.A1(_04218_),
    .A2(_04220_),
    .B(_04145_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10068_ (.I(net66),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10069_ (.I(_04222_),
    .Z(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _10070_ (.A1(_04199_),
    .A2(_03871_),
    .B1(_04211_),
    .B2(_00688_),
    .C1(_00817_),
    .C2(net40),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10071_ (.I(_00982_),
    .Z(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10072_ (.I(_04225_),
    .Z(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10073_ (.A1(_04223_),
    .A2(_03752_),
    .B1(_04224_),
    .B2(_04226_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10074_ (.I(_00793_),
    .Z(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10075_ (.I(_04136_),
    .Z(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10076_ (.A1(net87),
    .A2(_02193_),
    .B(_04229_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10077_ (.A1(_04150_),
    .A2(_04169_),
    .B(_04230_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10078_ (.A1(_04217_),
    .A2(_04231_),
    .Z(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10079_ (.A1(_04228_),
    .A2(_04232_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10080_ (.A1(_04209_),
    .A2(_02955_),
    .B(_04233_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10081_ (.A1(_03737_),
    .A2(_04227_),
    .B1(_04234_),
    .B2(_03818_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10082_ (.I(_04235_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10083_ (.I(_00800_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10084_ (.A1(_02212_),
    .A2(_04008_),
    .B1(_04236_),
    .B2(_04237_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10085_ (.A1(_04212_),
    .A2(_04221_),
    .B1(_04238_),
    .B2(_04161_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10086_ (.A1(_02212_),
    .A2(_03788_),
    .B1(_04239_),
    .B2(_04163_),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10087_ (.A1(net40),
    .A2(_04067_),
    .B(_04165_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10088_ (.A1(_04068_),
    .A2(_04240_),
    .B(_04241_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10089_ (.I(\as2650.addr_buff[3] ),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10090_ (.A1(_04242_),
    .A2(_04203_),
    .Z(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10091_ (.A1(_04242_),
    .A2(_04206_),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10092_ (.A1(_04129_),
    .A2(_04243_),
    .B1(_04244_),
    .B2(_04024_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10093_ (.A1(_04209_),
    .A2(_04210_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10094_ (.A1(net41),
    .A2(_04246_),
    .Z(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10095_ (.A1(_00719_),
    .A2(_04245_),
    .B1(_04247_),
    .B2(_03995_),
    .C(_03777_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10096_ (.A1(net67),
    .A2(_01608_),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10097_ (.A1(_02211_),
    .A2(_04229_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10098_ (.A1(_04250_),
    .A2(_04218_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10099_ (.A1(_04249_),
    .A2(_04251_),
    .Z(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10100_ (.A1(_03789_),
    .A2(_04252_),
    .B(_04145_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10101_ (.A1(_04009_),
    .A2(_04247_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10102_ (.I(\as2650.addr_buff[3] ),
    .Z(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10103_ (.I(net41),
    .Z(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10104_ (.A1(_04255_),
    .A2(_04103_),
    .B1(_04104_),
    .B2(_04256_),
    .C(_01291_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10105_ (.A1(_04254_),
    .A2(_04257_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10106_ (.A1(_02218_),
    .A2(_04101_),
    .B(_04258_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10107_ (.A1(_04217_),
    .A2(_04231_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10108_ (.A1(_04250_),
    .A2(_04260_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10109_ (.A1(_04249_),
    .A2(_04261_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10110_ (.A1(_03867_),
    .A2(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10111_ (.A1(_04256_),
    .A2(_04099_),
    .B(_03727_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10112_ (.A1(_04109_),
    .A2(_04259_),
    .B1(_04263_),
    .B2(_04264_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10113_ (.A1(_02218_),
    .A2(_04111_),
    .B1(_04265_),
    .B2(_03830_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10114_ (.A1(_04248_),
    .A2(_04253_),
    .B(_04266_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10115_ (.A1(_02218_),
    .A2(_03788_),
    .B1(_04267_),
    .B2(_04163_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10116_ (.A1(_04256_),
    .A2(_04067_),
    .B(_04165_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10117_ (.A1(_03721_),
    .A2(_04268_),
    .B(_04269_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10118_ (.I(\as2650.addr_buff[4] ),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10119_ (.A1(_04255_),
    .A2(_04118_),
    .A3(_04120_),
    .A4(_04202_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10120_ (.A1(_04270_),
    .A2(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10121_ (.A1(\as2650.addr_buff[3] ),
    .A2(_04124_),
    .A3(_04126_),
    .A4(_04202_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10122_ (.A1(_04270_),
    .A2(_04273_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10123_ (.I(_03991_),
    .Z(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10124_ (.A1(_03769_),
    .A2(_04272_),
    .B1(_04274_),
    .B2(_04275_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10125_ (.A1(_04256_),
    .A2(_04246_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10126_ (.A1(net92),
    .A2(_04277_),
    .Z(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10127_ (.A1(_03759_),
    .A2(_04276_),
    .B1(_04278_),
    .B2(_03772_),
    .C(_03774_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10128_ (.A1(_04216_),
    .A2(_04249_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10129_ (.A1(_02216_),
    .A2(_01609_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10130_ (.A1(_04250_),
    .A2(_04230_),
    .A3(_04281_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10131_ (.A1(_04215_),
    .A2(_04280_),
    .B(_04282_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10132_ (.A1(net68),
    .A2(_02940_),
    .Z(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10133_ (.A1(_04283_),
    .A2(_04284_),
    .Z(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10134_ (.A1(_04004_),
    .A2(_04285_),
    .B(_03781_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10135_ (.A1(_04279_),
    .A2(_04286_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10136_ (.A1(_04270_),
    .A2(_04103_),
    .B1(_04104_),
    .B2(net92),
    .C(_01291_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10137_ (.A1(_04102_),
    .A2(_04278_),
    .B(_04288_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10138_ (.A1(_02225_),
    .A2(_04101_),
    .B(_04289_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10139_ (.A1(_04150_),
    .A2(_04168_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10140_ (.A1(_04291_),
    .A2(_04280_),
    .B(_04282_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10141_ (.A1(_04284_),
    .A2(_04292_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10142_ (.A1(_00810_),
    .A2(_04293_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10143_ (.A1(net92),
    .A2(_04099_),
    .B(_03728_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10144_ (.A1(_00673_),
    .A2(_04290_),
    .B1(_04294_),
    .B2(_04295_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10145_ (.A1(_02225_),
    .A2(_04111_),
    .B1(_04296_),
    .B2(_00452_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10146_ (.I(_03779_),
    .Z(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10147_ (.A1(_04287_),
    .A2(_04297_),
    .B(_04298_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10148_ (.A1(_02225_),
    .A2(_04069_),
    .B(_04299_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10149_ (.I(_00678_),
    .Z(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10150_ (.A1(net92),
    .A2(_04067_),
    .B(_04301_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10151_ (.A1(_03721_),
    .A2(_04300_),
    .B(_04302_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10152_ (.A1(_02549_),
    .A2(_02578_),
    .A3(_03696_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10153_ (.A1(_02586_),
    .A2(_04303_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10154_ (.A1(_03699_),
    .A2(_04304_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10155_ (.A1(_03687_),
    .A2(_03690_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10156_ (.A1(_00906_),
    .A2(_00986_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10157_ (.A1(_03685_),
    .A2(_04307_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10158_ (.A1(_00631_),
    .A2(_00905_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10159_ (.A1(_04077_),
    .A2(_04309_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10160_ (.A1(_02552_),
    .A2(_00555_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10161_ (.A1(_00546_),
    .A2(_04311_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10162_ (.A1(_00782_),
    .A2(_02737_),
    .A3(_03678_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10163_ (.A1(_00808_),
    .A2(_00608_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10164_ (.A1(_00938_),
    .A2(_02333_),
    .A3(_04314_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10165_ (.A1(_04313_),
    .A2(_04315_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10166_ (.A1(_03870_),
    .A2(_00812_),
    .A3(_03651_),
    .A4(_04311_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10167_ (.A1(_00891_),
    .A2(_04317_),
    .B(_03598_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10168_ (.A1(_00556_),
    .A2(_00715_),
    .A3(_03650_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10169_ (.A1(_00546_),
    .A2(_02599_),
    .A3(_04319_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10170_ (.A1(_03677_),
    .A2(_04316_),
    .A3(_04318_),
    .A4(_04320_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10171_ (.A1(_00723_),
    .A2(_04308_),
    .B1(_04310_),
    .B2(_04312_),
    .C(_04321_),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _10172_ (.A1(_02561_),
    .A2(_02563_),
    .A3(_02594_),
    .A4(_03695_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10173_ (.A1(_04306_),
    .A2(_04322_),
    .A3(_04323_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10174_ (.A1(_03684_),
    .A2(_03715_),
    .A3(_04305_),
    .A4(_04324_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10175_ (.I(_02608_),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10176_ (.I(_04326_),
    .Z(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10177_ (.A1(net82),
    .A2(_04327_),
    .A3(_02811_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10178_ (.A1(_02352_),
    .A2(_00899_),
    .B(_04328_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10179_ (.A1(net28),
    .A2(_00611_),
    .B(_03646_),
    .C(_03781_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10180_ (.I(_00578_),
    .Z(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10181_ (.I(_04331_),
    .Z(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10182_ (.I(_04332_),
    .Z(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10183_ (.A1(net28),
    .A2(_04333_),
    .A3(_03968_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10184_ (.A1(_00801_),
    .A2(_04329_),
    .B(_04330_),
    .C(_04334_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10185_ (.A1(_02893_),
    .A2(_04325_),
    .B1(_04335_),
    .B2(_00507_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10186_ (.A1(net83),
    .A2(_04325_),
    .B(_04336_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10187_ (.I(net91),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10188_ (.A1(_00563_),
    .A2(_02547_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10189_ (.A1(_00560_),
    .A2(_00565_),
    .A3(_04338_),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10190_ (.A1(_00863_),
    .A2(_02722_),
    .A3(_00627_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10191_ (.A1(_00734_),
    .A2(_00450_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10192_ (.A1(_00601_),
    .A2(_04341_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10193_ (.I(_04341_),
    .Z(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10194_ (.A1(_00778_),
    .A2(_02008_),
    .A3(_04343_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10195_ (.A1(_00753_),
    .A2(_04340_),
    .A3(_04342_),
    .B1(_04344_),
    .B2(_00473_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10196_ (.A1(_04339_),
    .A2(_04345_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10197_ (.A1(_00548_),
    .A2(\as2650.cycle[12] ),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10198_ (.I(_03875_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10199_ (.I(_02572_),
    .Z(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10200_ (.A1(_00548_),
    .A2(\as2650.cycle[7] ),
    .B(_00525_),
    .C(_04349_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10201_ (.A1(_04347_),
    .A2(_00740_),
    .A3(_04348_),
    .A4(_04350_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10202_ (.A1(_03710_),
    .A2(_03697_),
    .A3(_04346_),
    .A4(_04351_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10203_ (.A1(_00519_),
    .A2(_03713_),
    .A3(_02759_),
    .A4(_04349_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10204_ (.A1(_03688_),
    .A2(_03714_),
    .A3(_03704_),
    .A4(_04353_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10205_ (.A1(_00580_),
    .A2(_04347_),
    .A3(_04338_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10206_ (.A1(_03692_),
    .A2(_02594_),
    .A3(_03676_),
    .A4(_04355_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10207_ (.A1(_03700_),
    .A2(_03716_),
    .A3(_04354_),
    .A4(_04356_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10208_ (.A1(_04352_),
    .A2(_04357_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10209_ (.A1(_03684_),
    .A2(_04358_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10210_ (.A1(net91),
    .A2(_00971_),
    .A3(_03649_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10211_ (.A1(_04331_),
    .A2(_00786_),
    .B(_04103_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10212_ (.A1(_03647_),
    .A2(_00700_),
    .B(_04361_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10213_ (.I(_00702_),
    .Z(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10214_ (.I(_04363_),
    .Z(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10215_ (.A1(net91),
    .A2(_04362_),
    .B(_04364_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10216_ (.A1(_04314_),
    .A2(_04365_),
    .B(_03755_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10217_ (.A1(net91),
    .A2(_02808_),
    .A3(_00496_),
    .A4(_00787_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10218_ (.A1(_00789_),
    .A2(_04367_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10219_ (.A1(_04366_),
    .A2(_04368_),
    .B(_04349_),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10220_ (.A1(_00707_),
    .A2(_00736_),
    .B1(_04360_),
    .B2(_04369_),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10221_ (.A1(_03977_),
    .A2(_04359_),
    .A3(_04370_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10222_ (.A1(_04337_),
    .A2(_04359_),
    .B(_04371_),
    .C(_03786_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10223_ (.A1(_00565_),
    .A2(_00700_),
    .B(_00741_),
    .C(_04348_),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10224_ (.A1(_03686_),
    .A2(_04309_),
    .B(_03649_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10225_ (.I(_00702_),
    .Z(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10226_ (.A1(_00880_),
    .A2(_03650_),
    .A3(_01131_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10227_ (.I(_03750_),
    .Z(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10228_ (.A1(_04376_),
    .A2(_00450_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10229_ (.A1(_04377_),
    .A2(_02333_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10230_ (.A1(_02806_),
    .A2(_02747_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10231_ (.A1(_00564_),
    .A2(_00556_),
    .B(_04379_),
    .C(_03644_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10232_ (.A1(_03877_),
    .A2(_00758_),
    .A3(_00926_),
    .A4(_02760_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10233_ (.A1(_03655_),
    .A2(_04378_),
    .A3(_04380_),
    .A4(_04381_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10234_ (.A1(_04374_),
    .A2(_00901_),
    .A3(_04375_),
    .A4(_04382_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10235_ (.A1(_04372_),
    .A2(_04373_),
    .A3(_04383_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10236_ (.I(_04384_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10237_ (.I0(_02845_),
    .I1(_04157_),
    .S(_04385_),
    .Z(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10238_ (.I(_04386_),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10239_ (.I(_04385_),
    .Z(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10240_ (.I(_04385_),
    .Z(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10241_ (.A1(_04186_),
    .A2(_04388_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10242_ (.A1(_03797_),
    .A2(_04387_),
    .B(_04389_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10243_ (.A1(_04200_),
    .A2(_04388_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10244_ (.A1(_01274_),
    .A2(_04387_),
    .B(_04390_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10245_ (.I(_04255_),
    .Z(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10246_ (.I(_04384_),
    .Z(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10247_ (.A1(_04391_),
    .A2(_04392_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10248_ (.A1(_03150_),
    .A2(_04387_),
    .B(_04393_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10249_ (.I(_03165_),
    .Z(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10250_ (.I(\as2650.addr_buff[4] ),
    .Z(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10251_ (.A1(_04395_),
    .A2(_04392_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10252_ (.A1(_04394_),
    .A2(_04387_),
    .B(_04396_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10253_ (.I(_02933_),
    .Z(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10254_ (.A1(_00978_),
    .A2(_04392_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10255_ (.A1(_04397_),
    .A2(_04388_),
    .B(_04398_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10256_ (.I(_02861_),
    .Z(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10257_ (.I(_00976_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10258_ (.I0(_04399_),
    .I1(_04400_),
    .S(_04385_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10259_ (.I(_04401_),
    .Z(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10260_ (.A1(_00639_),
    .A2(_04392_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10261_ (.A1(_00795_),
    .A2(_04388_),
    .B(_04402_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10262_ (.A1(\as2650.last_intr ),
    .A2(_02606_),
    .B(_04301_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10263_ (.A1(_00568_),
    .A2(_02606_),
    .B(_04403_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10264_ (.I(_00695_),
    .Z(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10265_ (.I(_04404_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10266_ (.A1(_02778_),
    .A2(_01024_),
    .B(_03673_),
    .C(_04405_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10267_ (.A1(_03673_),
    .A2(_02741_),
    .B(_03692_),
    .ZN(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10268_ (.A1(_02569_),
    .A2(_02964_),
    .B(_04406_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10269_ (.A1(_03712_),
    .A2(_04320_),
    .A3(_04407_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10270_ (.I(_03991_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10271_ (.A1(_04409_),
    .A2(_03685_),
    .A3(_04307_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10272_ (.A1(_03685_),
    .A2(_04309_),
    .B(_03689_),
    .C(_03707_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10273_ (.A1(_03706_),
    .A2(_04408_),
    .A3(_04410_),
    .A4(_04411_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10274_ (.A1(_00978_),
    .A2(_00822_),
    .B(_04412_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10275_ (.A1(_01121_),
    .A2(_04412_),
    .B(_04413_),
    .C(_04405_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10276_ (.A1(_04400_),
    .A2(_00822_),
    .B(_04412_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10277_ (.A1(_01008_),
    .A2(_04412_),
    .B(_04414_),
    .C(_04405_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10278_ (.A1(_02865_),
    .A2(_02844_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10279_ (.A1(_01022_),
    .A2(_03877_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10280_ (.A1(_04415_),
    .A2(_04416_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10281_ (.I(_02772_),
    .Z(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10282_ (.I(_04418_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10283_ (.A1(_00941_),
    .A2(_01345_),
    .B(_00515_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10284_ (.A1(_00767_),
    .A2(_04420_),
    .B(_00765_),
    .C(_03749_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10285_ (.A1(_04419_),
    .A2(_04421_),
    .B(_00966_),
    .C(_00911_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10286_ (.I(_04422_),
    .Z(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10287_ (.I0(_04417_),
    .I1(_01061_),
    .S(_04423_),
    .Z(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10288_ (.I(_04424_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10289_ (.I(_04422_),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10290_ (.I(_04425_),
    .Z(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10291_ (.A1(_02332_),
    .A2(_02847_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10292_ (.I(_02349_),
    .Z(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10293_ (.A1(_01136_),
    .A2(_04428_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10294_ (.A1(_04427_),
    .A2(_04429_),
    .Z(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10295_ (.A1(\as2650.holding_reg[1] ),
    .A2(_04426_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10296_ (.A1(_04426_),
    .A2(_04430_),
    .B(_04431_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10297_ (.I(_03877_),
    .Z(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10298_ (.A1(_01262_),
    .A2(_04432_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10299_ (.A1(_02618_),
    .A2(_02850_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10300_ (.A1(_04433_),
    .A2(_04434_),
    .Z(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10301_ (.A1(\as2650.holding_reg[2] ),
    .A2(_04423_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10302_ (.A1(_04426_),
    .A2(_04435_),
    .B(_04436_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10303_ (.I(_02855_),
    .Z(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10304_ (.A1(_02332_),
    .A2(_04437_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10305_ (.I(_04428_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10306_ (.A1(_01905_),
    .A2(_04439_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10307_ (.A1(_04438_),
    .A2(_04440_),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10308_ (.A1(\as2650.holding_reg[3] ),
    .A2(_04423_),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10309_ (.A1(_04426_),
    .A2(_04441_),
    .B(_04442_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10310_ (.A1(_01927_),
    .A2(_04439_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10311_ (.A1(_04327_),
    .A2(_04394_),
    .B(_04443_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10312_ (.I0(_04444_),
    .I1(\as2650.holding_reg[4] ),
    .S(_04423_),
    .Z(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10313_ (.I(_04445_),
    .Z(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10314_ (.A1(_04428_),
    .A2(_04397_),
    .B(_02609_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10315_ (.I0(_04446_),
    .I1(_01478_),
    .S(_04425_),
    .Z(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10316_ (.I(_04447_),
    .Z(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10317_ (.A1(_05674_),
    .A2(_04399_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10318_ (.A1(_03609_),
    .A2(_02903_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10319_ (.A1(_04448_),
    .A2(_04449_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10320_ (.I0(_04450_),
    .I1(\as2650.holding_reg[6] ),
    .S(_04425_),
    .Z(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10321_ (.I(_04451_),
    .Z(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10322_ (.A1(_02903_),
    .A2(_00795_),
    .B(_02353_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10323_ (.I0(_04452_),
    .I1(\as2650.holding_reg[7] ),
    .S(_04425_),
    .Z(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10324_ (.I(_04453_),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10325_ (.I(_04376_),
    .Z(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10326_ (.A1(_04454_),
    .A2(_00783_),
    .A3(_00786_),
    .A4(_04340_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10327_ (.A1(_00736_),
    .A2(_04455_),
    .B(_00507_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10328_ (.I(_04456_),
    .Z(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10329_ (.I(_04456_),
    .Z(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10330_ (.A1(_00737_),
    .A2(_02845_),
    .B(_04343_),
    .C(_04458_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10331_ (.A1(_00826_),
    .A2(_04457_),
    .B(_04459_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10332_ (.I(_02847_),
    .Z(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10333_ (.A1(_00737_),
    .A2(_04460_),
    .B(_04343_),
    .C(_04458_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10334_ (.A1(_02342_),
    .A2(_04457_),
    .B(_04461_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10335_ (.I(_02850_),
    .Z(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10336_ (.I(_00750_),
    .Z(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10337_ (.A1(_04462_),
    .A2(_04463_),
    .B1(_04457_),
    .B2(_00781_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10338_ (.I(_04464_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10339_ (.A1(_04377_),
    .A2(_00887_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10340_ (.A1(_00737_),
    .A2(_02614_),
    .B1(_04343_),
    .B2(_04465_),
    .C(_04456_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10341_ (.A1(_00460_),
    .A2(_04457_),
    .B(_04466_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10342_ (.A1(_04399_),
    .A2(_04463_),
    .B1(_04458_),
    .B2(_00827_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10343_ (.I(_04467_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10344_ (.A1(_00811_),
    .A2(_00751_),
    .B1(_04458_),
    .B2(_00825_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10345_ (.I(_04468_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10346_ (.I(_03692_),
    .Z(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10347_ (.I(_04469_),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10348_ (.I(_04406_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10349_ (.A1(_00670_),
    .A2(_03673_),
    .A3(_02741_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10350_ (.A1(_04471_),
    .A2(_04472_),
    .B(_00467_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10351_ (.A1(_00697_),
    .A2(_04470_),
    .A3(_04473_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10352_ (.A1(_00725_),
    .A2(_01004_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10353_ (.A1(_03991_),
    .A2(_04307_),
    .A3(_04474_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10354_ (.A1(_00715_),
    .A2(_00906_),
    .B(_04310_),
    .C(_04475_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10355_ (.A1(_00639_),
    .A2(_04375_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10356_ (.A1(_00881_),
    .A2(_00611_),
    .B(_04477_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10357_ (.A1(_04326_),
    .A2(_03637_),
    .B(_04380_),
    .C(_03659_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10358_ (.A1(_03649_),
    .A2(_04476_),
    .B(_04478_),
    .C(_04479_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10359_ (.I(_04480_),
    .Z(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10360_ (.A1(_00881_),
    .A2(_00979_),
    .Z(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10361_ (.I(_04482_),
    .Z(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10362_ (.I(_04482_),
    .Z(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10363_ (.A1(_01139_),
    .A2(_04484_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10364_ (.A1(_01101_),
    .A2(_04483_),
    .B(_04485_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10365_ (.I(_04480_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10366_ (.A1(net43),
    .A2(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10367_ (.A1(_04481_),
    .A2(_04486_),
    .B(_04488_),
    .C(_04405_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10368_ (.I(_04487_),
    .Z(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10369_ (.I(_04482_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10370_ (.I(_04482_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10371_ (.A1(_03138_),
    .A2(_04491_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10372_ (.A1(_03261_),
    .A2(_04490_),
    .B(_04492_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10373_ (.I(_04480_),
    .Z(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10374_ (.A1(net44),
    .A2(_04494_),
    .B(_04301_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10375_ (.A1(_04489_),
    .A2(_04493_),
    .B(_04495_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10376_ (.A1(_03148_),
    .A2(_04491_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10377_ (.A1(_03267_),
    .A2(_04490_),
    .B(_04496_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10378_ (.A1(net45),
    .A2(_04494_),
    .B(_04301_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10379_ (.A1(_04489_),
    .A2(_04497_),
    .B(_04498_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10380_ (.A1(_01431_),
    .A2(_04491_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10381_ (.A1(_03273_),
    .A2(_04490_),
    .B(_04499_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10382_ (.I(_00678_),
    .Z(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10383_ (.A1(net46),
    .A2(_04494_),
    .B(_04501_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10384_ (.A1(_04489_),
    .A2(_04500_),
    .B(_04502_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10385_ (.A1(_01460_),
    .A2(_04484_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10386_ (.A1(_03279_),
    .A2(_04483_),
    .B(_04503_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10387_ (.A1(net47),
    .A2(_04487_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10388_ (.I(_04404_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10389_ (.A1(_04481_),
    .A2(_04504_),
    .B(_04505_),
    .C(_04506_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10390_ (.A1(_02835_),
    .A2(_04491_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10391_ (.A1(_03285_),
    .A2(_04490_),
    .B(_04507_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10392_ (.A1(net21),
    .A2(_04494_),
    .B(_04501_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10393_ (.A1(_04489_),
    .A2(_04508_),
    .B(_04509_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10394_ (.A1(_02837_),
    .A2(_04484_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10395_ (.A1(_03609_),
    .A2(_04483_),
    .B(_04510_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10396_ (.A1(net22),
    .A2(_04487_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10397_ (.A1(_04481_),
    .A2(_04511_),
    .B(_04512_),
    .C(_04506_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10398_ (.A1(_02834_),
    .A2(_04484_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10399_ (.A1(_02347_),
    .A2(_04483_),
    .B(_04513_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10400_ (.A1(net23),
    .A2(_04480_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10401_ (.A1(_04481_),
    .A2(_04514_),
    .B(_04515_),
    .C(_04506_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10402_ (.A1(_02551_),
    .A2(_02556_),
    .A3(_03702_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10403_ (.A1(_02602_),
    .A2(_03712_),
    .A3(_03705_),
    .A4(_04516_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10404_ (.A1(_03714_),
    .A2(_04339_),
    .A3(_04355_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10405_ (.A1(_04351_),
    .A2(_04517_),
    .A3(_04518_),
    .Z(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10406_ (.I(_04411_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10407_ (.A1(_00519_),
    .A2(_00893_),
    .A3(_00565_),
    .A4(_04311_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10408_ (.A1(_00602_),
    .A2(_02573_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10409_ (.A1(_02732_),
    .A2(_00705_),
    .A3(_04521_),
    .B(_04522_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10410_ (.A1(_00662_),
    .A2(_00704_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10411_ (.A1(_00637_),
    .A2(_02013_),
    .A3(_04341_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10412_ (.A1(_02553_),
    .A2(_03598_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10413_ (.A1(_04524_),
    .A2(_04525_),
    .B(_04308_),
    .C(_04526_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10414_ (.A1(_04323_),
    .A2(_04520_),
    .A3(_04523_),
    .A4(_04527_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10415_ (.A1(_04305_),
    .A2(_04519_),
    .A3(_04528_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10416_ (.I(_04529_),
    .Z(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10417_ (.I(_04530_),
    .Z(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10418_ (.A1(_04469_),
    .A2(_03757_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10419_ (.I(_04532_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10420_ (.A1(_00799_),
    .A2(_02570_),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10421_ (.I(_04534_),
    .Z(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10422_ (.I(_01737_),
    .Z(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10423_ (.A1(\as2650.stack[7][0] ),
    .A2(_04536_),
    .B1(_01744_),
    .B2(\as2650.stack[6][0] ),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10424_ (.A1(\as2650.stack[5][0] ),
    .A2(_02784_),
    .B1(_02794_),
    .B2(\as2650.stack[4][0] ),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10425_ (.A1(_01786_),
    .A2(_04537_),
    .A3(_04538_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10426_ (.I(_02788_),
    .Z(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10427_ (.A1(\as2650.stack[1][0] ),
    .A2(_01789_),
    .B1(_01793_),
    .B2(\as2650.stack[0][0] ),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10428_ (.I(_01743_),
    .Z(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10429_ (.A1(\as2650.stack[3][0] ),
    .A2(_04536_),
    .B1(_04542_),
    .B2(\as2650.stack[2][0] ),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10430_ (.A1(_04540_),
    .A2(_04541_),
    .A3(_04543_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10431_ (.A1(_02779_),
    .A2(_04539_),
    .A3(_04544_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10432_ (.A1(\as2650.stack[9][0] ),
    .A2(_02784_),
    .B1(_02794_),
    .B2(\as2650.stack[8][0] ),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10433_ (.A1(\as2650.stack[11][0] ),
    .A2(_04536_),
    .B1(_01744_),
    .B2(\as2650.stack[10][0] ),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10434_ (.A1(_04540_),
    .A2(_04546_),
    .A3(_04547_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10435_ (.A1(\as2650.stack[15][0] ),
    .A2(_04536_),
    .B1(_04542_),
    .B2(\as2650.stack[14][0] ),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10436_ (.A1(\as2650.stack[13][0] ),
    .A2(_01789_),
    .B1(_01793_),
    .B2(\as2650.stack[12][0] ),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10437_ (.A1(_02906_),
    .A2(_04549_),
    .A3(_04550_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10438_ (.A1(_01775_),
    .A2(_04548_),
    .A3(_04551_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10439_ (.A1(_04545_),
    .A2(_04552_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10440_ (.I(_03665_),
    .Z(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10441_ (.A1(_03722_),
    .A2(_04076_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10442_ (.A1(_04076_),
    .A2(_03731_),
    .B(_04555_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10443_ (.A1(_03722_),
    .A2(_00779_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10444_ (.A1(_04376_),
    .A2(_04556_),
    .B(_04557_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10445_ (.A1(_04418_),
    .A2(_04558_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10446_ (.A1(_02037_),
    .A2(_00513_),
    .Z(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10447_ (.I0(_02038_),
    .I1(_04560_),
    .S(_00441_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10448_ (.I0(_02038_),
    .I1(_04560_),
    .S(_05703_),
    .Z(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10449_ (.A1(_00879_),
    .A2(_00827_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10450_ (.I0(_04561_),
    .I1(_04562_),
    .S(_04563_),
    .Z(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10451_ (.A1(_03739_),
    .A2(_00687_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10452_ (.A1(_03745_),
    .A2(_04565_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10453_ (.A1(_00520_),
    .A2(_04566_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10454_ (.A1(_04156_),
    .A2(_00520_),
    .A3(_00894_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10455_ (.A1(_04428_),
    .A2(_04564_),
    .B1(_04567_),
    .B2(_04568_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10456_ (.I(_04225_),
    .Z(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10457_ (.A1(_05777_),
    .A2(_00687_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10458_ (.A1(_03739_),
    .A2(_04571_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10459_ (.A1(_03739_),
    .A2(_04571_),
    .B(_04572_),
    .C(_04225_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10460_ (.A1(_03723_),
    .A2(_04570_),
    .B(_04573_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10461_ (.A1(_04559_),
    .A2(_04569_),
    .B1(_04574_),
    .B2(_04332_),
    .C(_04363_),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10462_ (.A1(_03749_),
    .A2(_04556_),
    .B(_03738_),
    .C(_00672_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10463_ (.A1(_04554_),
    .A2(_04575_),
    .A3(_04576_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10464_ (.A1(_03726_),
    .A2(_04535_),
    .B1(_02758_),
    .B2(_04553_),
    .C(_04577_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10465_ (.A1(_03916_),
    .A2(_04578_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10466_ (.A1(_03726_),
    .A2(_04533_),
    .B(_04530_),
    .C(_04579_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10467_ (.A1(_03726_),
    .A2(_04531_),
    .B(_04580_),
    .C(_04506_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10468_ (.A1(_02056_),
    .A2(_03722_),
    .Z(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10469_ (.I(_04581_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10470_ (.I(_00800_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10471_ (.I(_00783_),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10472_ (.A1(_04186_),
    .A2(_03873_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10473_ (.I(_00698_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10474_ (.I(_04586_),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10475_ (.I(_03746_),
    .Z(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10476_ (.A1(_02846_),
    .A2(_04587_),
    .B(_04588_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10477_ (.I(_04376_),
    .Z(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10478_ (.A1(_03787_),
    .A2(_03866_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10479_ (.A1(_00809_),
    .A2(_03821_),
    .B(_04591_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10480_ (.A1(_00780_),
    .A2(_04581_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10481_ (.A1(_04590_),
    .A2(_04592_),
    .B(_04593_),
    .C(_02334_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10482_ (.I(_00443_),
    .Z(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10483_ (.I(_04595_),
    .Z(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10484_ (.A1(net90),
    .A2(\as2650.ins_reg[2] ),
    .B(net56),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10485_ (.A1(_02057_),
    .A2(_02039_),
    .A3(_00804_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10486_ (.A1(_04597_),
    .A2(_04598_),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10487_ (.A1(_00445_),
    .A2(_04599_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10488_ (.A1(_04596_),
    .A2(_04582_),
    .B(_04600_),
    .C(_04432_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10489_ (.A1(_04585_),
    .A2(_04589_),
    .B(_04594_),
    .C(_04601_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10490_ (.A1(_04584_),
    .A2(_04602_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10491_ (.I(_02824_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10492_ (.A1(_04604_),
    .A2(_04581_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10493_ (.I(_04374_),
    .Z(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10494_ (.A1(_04327_),
    .A2(_04592_),
    .B(_04605_),
    .C(_04606_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10495_ (.I(_03745_),
    .Z(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10496_ (.I(_04608_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10497_ (.I(_04608_),
    .Z(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10498_ (.A1(net8),
    .A2(_05777_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10499_ (.A1(_03795_),
    .A2(_05782_),
    .Z(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10500_ (.A1(_04611_),
    .A2(_04612_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10501_ (.A1(_04611_),
    .A2(_04612_),
    .Z(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10502_ (.A1(_00689_),
    .A2(_04613_),
    .A3(_04614_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10503_ (.A1(_02846_),
    .A2(_04586_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10504_ (.A1(_04610_),
    .A2(_04615_),
    .A3(_04616_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10505_ (.A1(_04609_),
    .A2(_04582_),
    .B(_04617_),
    .C(_04333_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10506_ (.A1(_04583_),
    .A2(_04603_),
    .A3(_04607_),
    .A4(_04618_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10507_ (.I(_04534_),
    .Z(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10508_ (.A1(_00929_),
    .A2(_02727_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10509_ (.I(_04621_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10510_ (.A1(\as2650.stack[7][1] ),
    .A2(_01835_),
    .B1(_01790_),
    .B2(\as2650.stack[5][1] ),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10511_ (.A1(\as2650.stack[6][1] ),
    .A2(_01823_),
    .B1(_01794_),
    .B2(\as2650.stack[4][1] ),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10512_ (.A1(_02907_),
    .A2(_04623_),
    .A3(_04624_),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10513_ (.I(_04540_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10514_ (.A1(\as2650.stack[1][1] ),
    .A2(_01829_),
    .B1(_01826_),
    .B2(\as2650.stack[0][1] ),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10515_ (.A1(\as2650.stack[3][1] ),
    .A2(_01835_),
    .B1(_02909_),
    .B2(\as2650.stack[2][1] ),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10516_ (.A1(_04626_),
    .A2(_04627_),
    .A3(_04628_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10517_ (.A1(_02780_),
    .A2(_04625_),
    .A3(_04629_),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10518_ (.A1(\as2650.stack[9][1] ),
    .A2(_01829_),
    .B1(_01826_),
    .B2(\as2650.stack[8][1] ),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10519_ (.A1(\as2650.stack[11][1] ),
    .A2(_01835_),
    .B1(_01823_),
    .B2(\as2650.stack[10][1] ),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10520_ (.A1(_04626_),
    .A2(_04631_),
    .A3(_04632_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10521_ (.A1(\as2650.stack[15][1] ),
    .A2(_01810_),
    .B1(_01823_),
    .B2(\as2650.stack[14][1] ),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10522_ (.A1(\as2650.stack[13][1] ),
    .A2(_01829_),
    .B1(_01826_),
    .B2(\as2650.stack[12][1] ),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10523_ (.A1(_01765_),
    .A2(_04634_),
    .A3(_04635_),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10524_ (.A1(_01845_),
    .A2(_04633_),
    .A3(_04636_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10525_ (.A1(_04630_),
    .A2(_04637_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10526_ (.A1(_04622_),
    .A2(_04638_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10527_ (.I(_03915_),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10528_ (.A1(_04620_),
    .A2(_04581_),
    .B(_04639_),
    .C(_04640_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10529_ (.I(_04529_),
    .Z(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10530_ (.I(_04642_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10531_ (.A1(_04533_),
    .A2(_04582_),
    .B1(_04619_),
    .B2(_04641_),
    .C(_04643_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10532_ (.I(_04404_),
    .Z(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10533_ (.A1(_02057_),
    .A2(_04531_),
    .B(_04644_),
    .C(_04645_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10534_ (.A1(_03876_),
    .A2(_02055_),
    .A3(_02038_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10535_ (.A1(_02057_),
    .A2(_02039_),
    .B(_02070_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10536_ (.A1(_04646_),
    .A2(_04647_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10537_ (.I(_04648_),
    .Z(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10538_ (.I(_04649_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10539_ (.I(_02350_),
    .Z(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10540_ (.I(_04651_),
    .Z(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10541_ (.A1(_02069_),
    .A2(_04597_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10542_ (.I(_04595_),
    .Z(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10543_ (.A1(_02071_),
    .A2(_04597_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10544_ (.A1(_04654_),
    .A2(_04655_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10545_ (.A1(_00446_),
    .A2(_04649_),
    .B1(_04653_),
    .B2(_04656_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10546_ (.A1(_02851_),
    .A2(_04587_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10547_ (.A1(_04200_),
    .A2(_03960_),
    .B(_04588_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10548_ (.A1(_03876_),
    .A2(_03866_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10549_ (.A1(_04077_),
    .A2(_03865_),
    .B(_04660_),
    .ZN(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10550_ (.A1(_00780_),
    .A2(_04648_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10551_ (.A1(_04590_),
    .A2(_04661_),
    .B(_04662_),
    .C(_02334_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10552_ (.A1(_04658_),
    .A2(_04659_),
    .B(_04663_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10553_ (.A1(_04652_),
    .A2(_04657_),
    .B(_04664_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10554_ (.A1(_04432_),
    .A2(_04661_),
    .B(_04374_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10555_ (.A1(_02902_),
    .A2(_04649_),
    .B(_04666_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10556_ (.I(_04570_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10557_ (.A1(net10),
    .A2(_05754_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10558_ (.A1(_01271_),
    .A2(_05754_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10559_ (.A1(_03790_),
    .A2(_05782_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10560_ (.A1(_04669_),
    .A2(_04670_),
    .B(_04671_),
    .C(_04614_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10561_ (.A1(_04671_),
    .A2(_04614_),
    .B(_04669_),
    .C(_04670_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10562_ (.A1(_00895_),
    .A2(_04673_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10563_ (.A1(_04672_),
    .A2(_04674_),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10564_ (.A1(_01274_),
    .A2(_03744_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10565_ (.A1(_04226_),
    .A2(_04676_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10566_ (.A1(_04668_),
    .A2(_04648_),
    .B1(_04675_),
    .B2(_04677_),
    .C(_00521_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10567_ (.A1(_04667_),
    .A2(_04678_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10568_ (.A1(_00517_),
    .A2(_04665_),
    .B(_04679_),
    .C(_04583_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10569_ (.I(_01744_),
    .Z(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10570_ (.A1(\as2650.stack[7][2] ),
    .A2(_02799_),
    .B1(_04681_),
    .B2(\as2650.stack[6][2] ),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10571_ (.A1(\as2650.stack[5][2] ),
    .A2(_02913_),
    .B1(_02914_),
    .B2(\as2650.stack[4][2] ),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10572_ (.A1(_01787_),
    .A2(_04682_),
    .A3(_04683_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10573_ (.A1(\as2650.stack[3][2] ),
    .A2(_02908_),
    .B1(_02785_),
    .B2(\as2650.stack[1][2] ),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10574_ (.A1(\as2650.stack[2][2] ),
    .A2(_04681_),
    .B1(_02914_),
    .B2(\as2650.stack[0][2] ),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10575_ (.A1(_02789_),
    .A2(_04685_),
    .A3(_04686_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10576_ (.A1(_02780_),
    .A2(_04684_),
    .A3(_04687_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10577_ (.A1(\as2650.stack[9][2] ),
    .A2(_01790_),
    .B1(_01794_),
    .B2(\as2650.stack[8][2] ),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10578_ (.A1(\as2650.stack[11][2] ),
    .A2(_02908_),
    .B1(_04681_),
    .B2(\as2650.stack[10][2] ),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10579_ (.A1(_04626_),
    .A2(_04689_),
    .A3(_04690_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10580_ (.A1(\as2650.stack[14][2] ),
    .A2(_04681_),
    .B1(_02914_),
    .B2(\as2650.stack[12][2] ),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10581_ (.A1(\as2650.stack[15][2] ),
    .A2(_02908_),
    .B1(_02913_),
    .B2(\as2650.stack[13][2] ),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10582_ (.A1(_01787_),
    .A2(_04692_),
    .A3(_04693_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10583_ (.A1(_01776_),
    .A2(_04691_),
    .A3(_04694_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10584_ (.A1(_04688_),
    .A2(_04695_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10585_ (.A1(_04622_),
    .A2(_04696_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10586_ (.A1(_04620_),
    .A2(_04649_),
    .B(_04697_),
    .C(_04640_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10587_ (.A1(_04533_),
    .A2(_04650_),
    .B1(_04680_),
    .B2(_04698_),
    .C(_04643_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10588_ (.A1(_02071_),
    .A2(_04531_),
    .B(_04699_),
    .C(_04645_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10589_ (.I(_04642_),
    .Z(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10590_ (.I(_04700_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10591_ (.A1(_02081_),
    .A2(_04646_),
    .Z(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10592_ (.A1(_03914_),
    .A2(_04646_),
    .Z(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10593_ (.A1(_03914_),
    .A2(_04653_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10594_ (.A1(_02070_),
    .A2(_04597_),
    .B(_02082_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10595_ (.A1(_04596_),
    .A2(_04704_),
    .A3(_04705_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10596_ (.A1(_00446_),
    .A2(_04703_),
    .B(_04706_),
    .C(_04604_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10597_ (.I(_03750_),
    .Z(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10598_ (.I(_04708_),
    .Z(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10599_ (.A1(_03921_),
    .A2(_03920_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10600_ (.A1(_03914_),
    .A2(_03734_),
    .B(_04710_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10601_ (.A1(_04454_),
    .A2(_04702_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10602_ (.A1(_04709_),
    .A2(_04711_),
    .B(_04712_),
    .C(_04419_),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10603_ (.A1(_04391_),
    .A2(_04587_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10604_ (.A1(_03150_),
    .A2(_00896_),
    .B(_04610_),
    .C(_04714_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10605_ (.A1(_04584_),
    .A2(_04707_),
    .A3(_04713_),
    .A4(_04715_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10606_ (.A1(_05673_),
    .A2(_04711_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10607_ (.A1(_02619_),
    .A2(_04702_),
    .B(_04717_),
    .C(_04606_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10608_ (.A1(net11),
    .A2(_05767_),
    .Z(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10609_ (.A1(_04669_),
    .A2(_04673_),
    .A3(_04719_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10610_ (.A1(_04669_),
    .A2(_04673_),
    .B(_04719_),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10611_ (.A1(_03960_),
    .A2(_04721_),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10612_ (.I(_00894_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10613_ (.A1(_02855_),
    .A2(_04723_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10614_ (.I(_03746_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10615_ (.A1(_04720_),
    .A2(_04722_),
    .B(_04724_),
    .C(_04725_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10616_ (.A1(_04609_),
    .A2(_04702_),
    .B(_04726_),
    .C(_04333_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10617_ (.A1(_04583_),
    .A2(_04716_),
    .A3(_04718_),
    .A4(_04727_),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10618_ (.A1(\as2650.stack[7][3] ),
    .A2(_01839_),
    .B1(_01752_),
    .B2(\as2650.stack[5][3] ),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10619_ (.A1(\as2650.stack[6][3] ),
    .A2(_01781_),
    .B1(_01757_),
    .B2(\as2650.stack[4][3] ),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10620_ (.A1(_01734_),
    .A2(_04729_),
    .A3(_04730_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10621_ (.A1(\as2650.stack[1][3] ),
    .A2(_01815_),
    .B1(_01818_),
    .B2(\as2650.stack[0][3] ),
    .C1(\as2650.stack[2][3] ),
    .C2(_01876_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10622_ (.A1(\as2650.stack[3][3] ),
    .A2(_01839_),
    .B(_02907_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10623_ (.A1(_04732_),
    .A2(_04733_),
    .B(_01776_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10624_ (.A1(\as2650.stack[9][3] ),
    .A2(_01815_),
    .B1(_01818_),
    .B2(\as2650.stack[8][3] ),
    .C1(\as2650.stack[10][3] ),
    .C2(_01876_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10625_ (.A1(\as2650.stack[11][3] ),
    .A2(_01839_),
    .B(_02907_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10626_ (.A1(\as2650.stack[15][3] ),
    .A2(_02782_),
    .B1(_01780_),
    .B2(\as2650.stack[14][3] ),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10627_ (.A1(\as2650.stack[13][3] ),
    .A2(_01751_),
    .B1(_02795_),
    .B2(\as2650.stack[12][3] ),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10628_ (.A1(_01733_),
    .A2(_04737_),
    .A3(_04738_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10629_ (.A1(_04735_),
    .A2(_04736_),
    .B(_04739_),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10630_ (.A1(_04731_),
    .A2(_04734_),
    .B1(_04740_),
    .B2(_01845_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10631_ (.I(_02758_),
    .Z(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10632_ (.A1(_04620_),
    .A2(_04703_),
    .B1(_04741_),
    .B2(_04742_),
    .C(_04640_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10633_ (.I(_04529_),
    .Z(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10634_ (.A1(_04533_),
    .A2(_04702_),
    .B1(_04728_),
    .B2(_04743_),
    .C(_04744_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10635_ (.A1(_02082_),
    .A2(_04701_),
    .B(_04745_),
    .C(_04645_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10636_ (.A1(net58),
    .A2(net57),
    .A3(net56),
    .A4(net55),
    .Z(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10637_ (.A1(_03958_),
    .A2(_04746_),
    .Z(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10638_ (.I(_04747_),
    .Z(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10639_ (.I(_04748_),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10640_ (.A1(_02093_),
    .A2(_04704_),
    .Z(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10641_ (.A1(_04596_),
    .A2(_04750_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10642_ (.I(_02824_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10643_ (.A1(_04654_),
    .A2(_04749_),
    .B(_04751_),
    .C(_04752_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10644_ (.A1(_03921_),
    .A2(_03964_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10645_ (.A1(_03958_),
    .A2(_02955_),
    .B(_04754_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10646_ (.A1(_04454_),
    .A2(_04747_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10647_ (.A1(_04709_),
    .A2(_04755_),
    .B(_04756_),
    .C(_04419_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10648_ (.A1(_04395_),
    .A2(_04587_),
    .ZN(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10649_ (.A1(_04394_),
    .A2(_00896_),
    .B(_04725_),
    .C(_04758_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10650_ (.A1(_04584_),
    .A2(_04753_),
    .A3(_04757_),
    .A4(_04759_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10651_ (.A1(_05673_),
    .A2(_04755_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10652_ (.A1(_02619_),
    .A2(_04748_),
    .B(_04761_),
    .C(_04606_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10653_ (.A1(_02852_),
    .A2(_05767_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10654_ (.A1(_01434_),
    .A2(_05761_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10655_ (.A1(_01434_),
    .A2(_05761_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10656_ (.A1(_04763_),
    .A2(_04721_),
    .B(_04764_),
    .C(_04765_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10657_ (.A1(_04764_),
    .A2(_04765_),
    .B(_04763_),
    .C(_04721_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10658_ (.A1(_03960_),
    .A2(_04767_),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10659_ (.A1(_02858_),
    .A2(_04009_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10660_ (.A1(_04766_),
    .A2(_04768_),
    .B(_04769_),
    .C(_04588_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10661_ (.I(_04332_),
    .Z(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10662_ (.A1(_04609_),
    .A2(_04748_),
    .B(_04770_),
    .C(_04771_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10663_ (.A1(_04583_),
    .A2(_04760_),
    .A3(_04762_),
    .A4(_04772_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10664_ (.A1(\as2650.stack[6][4] ),
    .A2(_01780_),
    .B1(_01751_),
    .B2(\as2650.stack[5][4] ),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10665_ (.A1(\as2650.stack[7][4] ),
    .A2(_01809_),
    .B1(_01756_),
    .B2(\as2650.stack[4][4] ),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10666_ (.A1(_01764_),
    .A2(_04774_),
    .A3(_04775_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10667_ (.A1(\as2650.stack[1][4] ),
    .A2(_01814_),
    .B1(_01817_),
    .B2(\as2650.stack[0][4] ),
    .C1(\as2650.stack[2][4] ),
    .C2(_01875_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10668_ (.A1(\as2650.stack[3][4] ),
    .A2(_01738_),
    .B(_01786_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10669_ (.A1(_04777_),
    .A2(_04778_),
    .B(_01775_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10670_ (.A1(\as2650.stack[9][4] ),
    .A2(_01814_),
    .B1(_01817_),
    .B2(\as2650.stack[8][4] ),
    .C1(\as2650.stack[10][4] ),
    .C2(_01875_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10671_ (.A1(\as2650.stack[11][4] ),
    .A2(_01738_),
    .B(_01786_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10672_ (.A1(\as2650.stack[15][4] ),
    .A2(_02781_),
    .B1(_01779_),
    .B2(\as2650.stack[14][4] ),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10673_ (.A1(\as2650.stack[13][4] ),
    .A2(_01750_),
    .B1(_01755_),
    .B2(\as2650.stack[12][4] ),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10674_ (.A1(_01732_),
    .A2(_04782_),
    .A3(_04783_),
    .Z(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10675_ (.A1(_04780_),
    .A2(_04781_),
    .B(_04784_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10676_ (.A1(_04776_),
    .A2(_04779_),
    .B1(_04785_),
    .B2(_01844_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10677_ (.A1(_04535_),
    .A2(_04749_),
    .B1(_04786_),
    .B2(_04742_),
    .C(_04640_),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10678_ (.A1(_04532_),
    .A2(_04748_),
    .B1(_04773_),
    .B2(_04787_),
    .C(_04744_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10679_ (.A1(_02094_),
    .A2(_04701_),
    .B(_04788_),
    .C(_04645_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10680_ (.I(_04530_),
    .Z(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10681_ (.I(_03661_),
    .Z(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10682_ (.A1(net60),
    .A2(_04746_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10683_ (.A1(_04007_),
    .A2(_04791_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10684_ (.I(_04792_),
    .Z(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10685_ (.I(_01291_),
    .Z(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10686_ (.A1(_01464_),
    .A2(_05737_),
    .Z(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10687_ (.A1(_04764_),
    .A2(_04766_),
    .A3(_04795_),
    .Z(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10688_ (.A1(_04764_),
    .A2(_04766_),
    .B(_04795_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10689_ (.A1(_04796_),
    .A2(_04797_),
    .B(_04586_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10690_ (.A1(_04397_),
    .A2(_00895_),
    .B(_04570_),
    .C(_04798_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10691_ (.A1(_04794_),
    .A2(_04793_),
    .B(_04799_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10692_ (.A1(_02105_),
    .A2(_03957_),
    .A3(_02080_),
    .A4(_04653_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10693_ (.I(_00444_),
    .Z(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10694_ (.A1(_02094_),
    .A2(_04704_),
    .B(_02107_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10695_ (.A1(_04802_),
    .A2(_04803_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10696_ (.I(_04792_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10697_ (.I(_00444_),
    .Z(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10698_ (.A1(_04801_),
    .A2(_04804_),
    .B1(_04805_),
    .B2(_04806_),
    .C(_02824_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10699_ (.I(_00779_),
    .Z(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10700_ (.A1(_02106_),
    .A2(_00628_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10701_ (.A1(_02952_),
    .A2(_04015_),
    .B(_04809_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10702_ (.I(_03750_),
    .Z(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10703_ (.A1(_04811_),
    .A2(_04792_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10704_ (.A1(_04808_),
    .A2(_04810_),
    .B(_04812_),
    .C(_04418_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10705_ (.A1(_00978_),
    .A2(_04586_),
    .B(_04105_),
    .ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10706_ (.A1(_04397_),
    .A2(_04723_),
    .B(_04814_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10707_ (.A1(_00521_),
    .A2(_04807_),
    .A3(_04813_),
    .A4(_04815_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10708_ (.A1(_00522_),
    .A2(_04800_),
    .B(_04816_),
    .C(_04109_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10709_ (.A1(_02351_),
    .A2(_04792_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10710_ (.I(_04363_),
    .Z(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10711_ (.A1(_03642_),
    .A2(_04810_),
    .B(_04818_),
    .C(_04819_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10712_ (.A1(_04237_),
    .A2(_04817_),
    .A3(_04820_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10713_ (.I(_01737_),
    .Z(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10714_ (.A1(\as2650.stack[7][5] ),
    .A2(_04822_),
    .B1(_01793_),
    .B2(\as2650.stack[4][5] ),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10715_ (.A1(\as2650.stack[6][5] ),
    .A2(_04542_),
    .B1(_01789_),
    .B2(\as2650.stack[5][5] ),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10716_ (.A1(_02906_),
    .A2(_04823_),
    .A3(_04824_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10717_ (.A1(\as2650.stack[3][5] ),
    .A2(_04822_),
    .B1(_01825_),
    .B2(\as2650.stack[0][5] ),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10718_ (.A1(\as2650.stack[2][5] ),
    .A2(_04542_),
    .B1(_01828_),
    .B2(\as2650.stack[1][5] ),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10719_ (.A1(_04540_),
    .A2(_04826_),
    .A3(_04827_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10720_ (.A1(_02779_),
    .A2(_04825_),
    .A3(_04828_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10721_ (.A1(\as2650.stack[9][5] ),
    .A2(_01828_),
    .B1(_01825_),
    .B2(\as2650.stack[8][5] ),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10722_ (.A1(\as2650.stack[11][5] ),
    .A2(_04822_),
    .B1(_01822_),
    .B2(\as2650.stack[10][5] ),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10723_ (.A1(_02789_),
    .A2(_04830_),
    .A3(_04831_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10724_ (.A1(\as2650.stack[15][5] ),
    .A2(_04822_),
    .B1(_01822_),
    .B2(\as2650.stack[14][5] ),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10725_ (.A1(\as2650.stack[13][5] ),
    .A2(_01828_),
    .B1(_01825_),
    .B2(\as2650.stack[12][5] ),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10726_ (.A1(_02906_),
    .A2(_04833_),
    .A3(_04834_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10727_ (.A1(_01844_),
    .A2(_04832_),
    .A3(_04835_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10728_ (.A1(_04829_),
    .A2(_04836_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10729_ (.A1(_04535_),
    .A2(_04793_),
    .B1(_04837_),
    .B2(_04742_),
    .C(_04062_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10730_ (.A1(_04821_),
    .A2(_04838_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10731_ (.A1(_04790_),
    .A2(_04793_),
    .B(_04839_),
    .C(_00732_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10732_ (.I(_02557_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10733_ (.A1(\as2650.ivec[0] ),
    .A2(_04470_),
    .B1(_04841_),
    .B2(_04793_),
    .C(_04530_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10734_ (.A1(_02107_),
    .A2(_04789_),
    .B1(_04840_),
    .B2(_04842_),
    .C(_00739_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10735_ (.A1(_04007_),
    .A2(_04791_),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10736_ (.A1(_02116_),
    .A2(_04843_),
    .Z(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10737_ (.I(_04844_),
    .Z(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10738_ (.I(_04844_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10739_ (.A1(_04229_),
    .A2(_05746_),
    .Z(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10740_ (.A1(_04229_),
    .A2(_05746_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10741_ (.A1(_01465_),
    .A2(_05737_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10742_ (.A1(_04847_),
    .A2(_04848_),
    .B(_04849_),
    .C(_04797_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10743_ (.A1(_04849_),
    .A2(_04797_),
    .B(_04847_),
    .C(_04848_),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10744_ (.A1(_00894_),
    .A2(_04851_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10745_ (.A1(_04025_),
    .A2(_04009_),
    .B1(_04850_),
    .B2(_04852_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10746_ (.I0(_04846_),
    .I1(_04853_),
    .S(_04608_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10747_ (.A1(_04023_),
    .A2(_04801_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10748_ (.A1(_04802_),
    .A2(_04855_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10749_ (.A1(_00445_),
    .A2(_04846_),
    .B(_04856_),
    .C(_02901_),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10750_ (.A1(_01697_),
    .A2(_04056_),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10751_ (.A1(_04023_),
    .A2(_03733_),
    .B(_04858_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10752_ (.A1(_04811_),
    .A2(_04844_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10753_ (.A1(_00780_),
    .A2(_04859_),
    .B(_04860_),
    .C(_04418_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10754_ (.A1(_04025_),
    .A2(_03744_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10755_ (.A1(_04400_),
    .A2(_00699_),
    .B(_04105_),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10756_ (.A1(_04862_),
    .A2(_04863_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10757_ (.A1(_00521_),
    .A2(_04857_),
    .A3(_04861_),
    .A4(_04864_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10758_ (.A1(_00522_),
    .A2(_04854_),
    .B(_04865_),
    .C(_03737_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10759_ (.A1(_02351_),
    .A2(_04845_),
    .ZN(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10760_ (.A1(_03642_),
    .A2(_04859_),
    .B(_04867_),
    .C(_04819_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10761_ (.A1(_04237_),
    .A2(_04866_),
    .A3(_04868_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10762_ (.A1(_04742_),
    .A2(_02804_),
    .B1(_04845_),
    .B2(_04534_),
    .C(_04062_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10763_ (.A1(_04869_),
    .A2(_04870_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10764_ (.A1(_04790_),
    .A2(_04845_),
    .B(_04871_),
    .C(_00732_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10765_ (.I(_04642_),
    .Z(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10766_ (.A1(\as2650.ivec[1] ),
    .A2(_04470_),
    .B1(_04841_),
    .B2(_04845_),
    .C(_04873_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10767_ (.A1(_02116_),
    .A2(_04789_),
    .B1(_04872_),
    .B2(_04874_),
    .C(_00739_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10768_ (.I(net63),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10769_ (.A1(_02115_),
    .A2(_04007_),
    .A3(_04791_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10770_ (.A1(_04875_),
    .A2(_04876_),
    .Z(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10771_ (.I(_04877_),
    .Z(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10772_ (.I(_00782_),
    .Z(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10773_ (.A1(_02115_),
    .A2(_04801_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10774_ (.A1(_02125_),
    .A2(_04880_),
    .Z(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10775_ (.A1(_02125_),
    .A2(_04880_),
    .B(_04802_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10776_ (.A1(_04881_),
    .A2(_04882_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10777_ (.I(_04877_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10778_ (.A1(_00445_),
    .A2(_04884_),
    .B(_03641_),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10779_ (.A1(_03870_),
    .A2(_00699_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10780_ (.A1(_03921_),
    .A2(_00895_),
    .B(_04608_),
    .C(_04886_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10781_ (.A1(_04875_),
    .A2(_00628_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10782_ (.A1(_02952_),
    .A2(_04097_),
    .B(_04888_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10783_ (.A1(_04811_),
    .A2(_04877_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10784_ (.I(_02772_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10785_ (.A1(_04808_),
    .A2(_04889_),
    .B(_04890_),
    .C(_04891_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10786_ (.A1(_04883_),
    .A2(_04885_),
    .B(_04887_),
    .C(_04892_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10787_ (.A1(_04879_),
    .A2(_04893_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10788_ (.A1(_04651_),
    .A2(_04878_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10789_ (.A1(_02902_),
    .A2(_04889_),
    .B(_04895_),
    .C(_04819_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10790_ (.I(_03746_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10791_ (.A1(net3),
    .A2(_05721_),
    .Z(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10792_ (.A1(_04847_),
    .A2(_04851_),
    .B(_04898_),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10793_ (.A1(_04847_),
    .A2(_04851_),
    .A3(_04898_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10794_ (.A1(_04899_),
    .A2(_04900_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10795_ (.A1(_03824_),
    .A2(_04901_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10796_ (.A1(_03820_),
    .A2(_00689_),
    .B(_04897_),
    .C(_04902_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10797_ (.I(_04331_),
    .Z(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10798_ (.A1(_04610_),
    .A2(_04884_),
    .B(_04903_),
    .C(_04904_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10799_ (.A1(_04237_),
    .A2(_04894_),
    .A3(_04896_),
    .A4(_04905_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10800_ (.A1(_02571_),
    .A2(_02924_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10801_ (.A1(_02621_),
    .A2(_04878_),
    .B(_04907_),
    .C(_04554_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10802_ (.A1(_02809_),
    .A2(_04906_),
    .A3(_04908_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10803_ (.A1(_04790_),
    .A2(_04878_),
    .B(_04909_),
    .C(_00732_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10804_ (.A1(\as2650.ivec[2] ),
    .A2(_04470_),
    .B1(_04841_),
    .B2(_04878_),
    .C(_04873_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10805_ (.I(_00711_),
    .Z(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10806_ (.A1(_04875_),
    .A2(_04789_),
    .B1(_04910_),
    .B2(_04911_),
    .C(_04912_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10807_ (.I(_02194_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10808_ (.A1(_04875_),
    .A2(_04876_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10809_ (.A1(_04913_),
    .A2(_04914_),
    .Z(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10810_ (.I(_04595_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10811_ (.A1(_02194_),
    .A2(_04881_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10812_ (.A1(_04916_),
    .A2(_04917_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10813_ (.A1(_04654_),
    .A2(_04915_),
    .B(_04918_),
    .C(_04651_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10814_ (.A1(_04913_),
    .A2(_04077_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10815_ (.A1(_00809_),
    .A2(_04152_),
    .B(_04920_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10816_ (.A1(_02194_),
    .A2(_04914_),
    .Z(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10817_ (.A1(_04808_),
    .A2(_04922_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10818_ (.A1(_04709_),
    .A2(_04921_),
    .B(_04923_),
    .C(_02334_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10819_ (.A1(_03740_),
    .A2(_04723_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10820_ (.A1(_04157_),
    .A2(_04102_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10821_ (.A1(_04725_),
    .A2(_04925_),
    .A3(_04926_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10822_ (.A1(_04879_),
    .A2(_04919_),
    .A3(_04924_),
    .A4(_04927_),
    .Z(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10823_ (.A1(_00627_),
    .A2(_05721_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10824_ (.A1(_04929_),
    .A2(_04899_),
    .B(_00698_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10825_ (.A1(_04116_),
    .A2(_04930_),
    .Z(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10826_ (.A1(_04668_),
    .A2(_04931_),
    .B(_04771_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10827_ (.A1(_04668_),
    .A2(_04915_),
    .B(_04932_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10828_ (.I(_04922_),
    .Z(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10829_ (.A1(_05673_),
    .A2(_04934_),
    .B(_04819_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10830_ (.A1(_02619_),
    .A2(_04921_),
    .B(_04935_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10831_ (.A1(_00452_),
    .A2(_04928_),
    .A3(_04933_),
    .A4(_04936_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10832_ (.A1(_03639_),
    .A2(_04934_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10833_ (.A1(_03639_),
    .A2(_01800_),
    .B(_04938_),
    .C(_00760_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10834_ (.A1(_04161_),
    .A2(_04934_),
    .B(_04939_),
    .C(_03780_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10835_ (.I(_02557_),
    .Z(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10836_ (.A1(\as2650.ivec[3] ),
    .A2(_04469_),
    .B1(_04941_),
    .B2(_04934_),
    .C(_04642_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10837_ (.A1(_04937_),
    .A2(_04940_),
    .B(_04942_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10838_ (.A1(_03972_),
    .A2(_04943_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10839_ (.A1(_04913_),
    .A2(_04531_),
    .B(_04944_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10840_ (.A1(_02193_),
    .A2(_04914_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10841_ (.A1(_04167_),
    .A2(_04945_),
    .Z(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10842_ (.I(_04946_),
    .Z(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10843_ (.I(_03665_),
    .Z(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10844_ (.A1(_02204_),
    .A2(net88),
    .A3(_04881_),
    .Z(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10845_ (.A1(_02195_),
    .A2(_04881_),
    .B(_02204_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10846_ (.A1(_04949_),
    .A2(_04950_),
    .B(_04806_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10847_ (.A1(_04916_),
    .A2(_04947_),
    .B(_04951_),
    .C(_04326_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10848_ (.A1(_04175_),
    .A2(_04723_),
    .B(_04616_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10849_ (.A1(_04588_),
    .A2(_04953_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10850_ (.A1(_00794_),
    .A2(_04192_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10851_ (.A1(_04167_),
    .A2(_04228_),
    .B(_04955_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10852_ (.I(_04946_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10853_ (.A1(_04708_),
    .A2(_04957_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10854_ (.A1(_04590_),
    .A2(_04956_),
    .B(_04958_),
    .C(_04891_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10855_ (.A1(_04952_),
    .A2(_04954_),
    .A3(_04959_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10856_ (.A1(_04116_),
    .A2(_04173_),
    .A3(_04930_),
    .Z(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10857_ (.A1(_04157_),
    .A2(_04930_),
    .B(_04186_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10858_ (.A1(_04226_),
    .A2(_04946_),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10859_ (.A1(_04794_),
    .A2(_04961_),
    .A3(_04962_),
    .B(_04963_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10860_ (.A1(_04326_),
    .A2(_04956_),
    .B(_04374_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10861_ (.A1(_04752_),
    .A2(_04957_),
    .B(_04965_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10862_ (.A1(_04879_),
    .A2(_04960_),
    .B1(_04964_),
    .B2(_04771_),
    .C(_04966_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10863_ (.I(_01847_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10864_ (.A1(_04968_),
    .A2(_02758_),
    .B1(_04947_),
    .B2(_04534_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10865_ (.A1(_04948_),
    .A2(_04967_),
    .B(_04969_),
    .C(_02809_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10866_ (.A1(_04790_),
    .A2(_04947_),
    .B(_04970_),
    .C(_04298_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10867_ (.I(_04469_),
    .Z(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10868_ (.A1(\as2650.ivec[4] ),
    .A2(_04972_),
    .B1(_04841_),
    .B2(_04947_),
    .C(_04873_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10869_ (.A1(_04167_),
    .A2(_04789_),
    .B1(_04971_),
    .B2(_04973_),
    .C(_04912_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10870_ (.A1(net65),
    .A2(net64),
    .A3(_04914_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10871_ (.A1(_04223_),
    .A2(_04974_),
    .Z(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10872_ (.A1(_04199_),
    .A2(_04102_),
    .B(_04676_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10873_ (.A1(_00794_),
    .A2(_04232_),
    .ZN(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10874_ (.A1(_04223_),
    .A2(_03733_),
    .B(_04977_),
    .ZN(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10875_ (.A1(_02211_),
    .A2(_04974_),
    .Z(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10876_ (.A1(_04708_),
    .A2(_04979_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10877_ (.A1(_04808_),
    .A2(_04978_),
    .B(_04980_),
    .C(_04891_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10878_ (.A1(_04222_),
    .A2(_04949_),
    .Z(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10879_ (.A1(_04806_),
    .A2(_04982_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10880_ (.A1(_04916_),
    .A2(_04975_),
    .B(_04983_),
    .C(_03641_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10881_ (.A1(_04794_),
    .A2(_04976_),
    .B(_04981_),
    .C(_04984_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10882_ (.A1(\as2650.addr_buff[0] ),
    .A2(\as2650.addr_buff[1] ),
    .A3(\as2650.addr_buff[2] ),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10883_ (.A1(_04929_),
    .A2(_04899_),
    .B(_00893_),
    .C(_04986_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10884_ (.I(_04987_),
    .Z(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10885_ (.A1(_04199_),
    .A2(_04961_),
    .B(_04897_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10886_ (.A1(_04725_),
    .A2(_04979_),
    .B1(_04988_),
    .B2(_04989_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10887_ (.A1(_03816_),
    .A2(_04978_),
    .B(_04363_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10888_ (.A1(_04752_),
    .A2(_04979_),
    .B(_04991_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10889_ (.A1(_04879_),
    .A2(_04985_),
    .B1(_04990_),
    .B2(_04771_),
    .C(_04992_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10890_ (.A1(_04948_),
    .A2(_04993_),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10891_ (.I(_04622_),
    .Z(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10892_ (.A1(_01884_),
    .A2(_04995_),
    .B1(_04979_),
    .B2(_03667_),
    .C(_00882_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10893_ (.A1(_03662_),
    .A2(_04975_),
    .B1(_04994_),
    .B2(_04996_),
    .C(_03832_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10894_ (.A1(\as2650.ivec[5] ),
    .A2(_04972_),
    .B1(_04941_),
    .B2(_04975_),
    .C(_04873_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10895_ (.A1(_04223_),
    .A2(_04700_),
    .B1(_04997_),
    .B2(_04998_),
    .C(_04912_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10896_ (.I(_02217_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10897_ (.A1(_04222_),
    .A2(_04974_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10898_ (.A1(_02217_),
    .A2(_05000_),
    .Z(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10899_ (.I(_05001_),
    .Z(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10900_ (.A1(_04999_),
    .A2(_00809_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10901_ (.A1(_03820_),
    .A2(_04262_),
    .B(_05003_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10902_ (.A1(_04454_),
    .A2(_05002_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10903_ (.A1(_04709_),
    .A2(_05004_),
    .B(_05005_),
    .C(_04419_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10904_ (.I(_05001_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10905_ (.A1(_02212_),
    .A2(_04949_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10906_ (.A1(_04999_),
    .A2(_05008_),
    .Z(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10907_ (.A1(_04596_),
    .A2(_05009_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10908_ (.A1(_04654_),
    .A2(_05007_),
    .B(_05010_),
    .C(_04752_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10909_ (.A1(_04391_),
    .A2(_03873_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10910_ (.A1(_04609_),
    .A2(_05012_),
    .A3(_04724_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10911_ (.A1(_05006_),
    .A2(_05011_),
    .A3(_05013_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10912_ (.A1(_04432_),
    .A2(_05002_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10913_ (.A1(_04604_),
    .A2(_05004_),
    .B(_05015_),
    .C(_04364_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10914_ (.A1(_04242_),
    .A2(_04987_),
    .B(_04570_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10915_ (.A1(_04391_),
    .A2(_04988_),
    .B(_05017_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10916_ (.A1(_04610_),
    .A2(_05007_),
    .B(_05018_),
    .C(_04904_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10917_ (.A1(_03755_),
    .A2(_05016_),
    .A3(_05019_),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10918_ (.A1(_04584_),
    .A2(_05014_),
    .B(_05020_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10919_ (.A1(_01904_),
    .A2(_04995_),
    .B1(_05007_),
    .B2(_03667_),
    .C(_00882_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10920_ (.A1(_03662_),
    .A2(_05002_),
    .B1(_05021_),
    .B2(_05022_),
    .C(_03832_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10921_ (.A1(\as2650.ivec[6] ),
    .A2(_04972_),
    .B1(_04941_),
    .B2(_05002_),
    .C(_04643_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10922_ (.A1(_04999_),
    .A2(_04700_),
    .B1(_05023_),
    .B2(_05024_),
    .C(_04912_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10923_ (.I(_02224_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10924_ (.I(_05025_),
    .Z(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10925_ (.A1(_02217_),
    .A2(_05000_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10926_ (.A1(_05026_),
    .A2(_05027_),
    .Z(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10927_ (.A1(_00794_),
    .A2(_04293_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10928_ (.A1(_05026_),
    .A2(_04228_),
    .B(_05029_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10929_ (.A1(_02224_),
    .A2(_02216_),
    .A3(_05000_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10930_ (.A1(_05026_),
    .A2(_05027_),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10931_ (.A1(_05031_),
    .A2(_05032_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10932_ (.A1(_04604_),
    .A2(_05033_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10933_ (.A1(_04327_),
    .A2(_05030_),
    .B(_05034_),
    .C(_04606_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10934_ (.A1(_04395_),
    .A2(_03824_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10935_ (.A1(_05036_),
    .A2(_04769_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10936_ (.A1(_04708_),
    .A2(_05033_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10937_ (.A1(_04590_),
    .A2(_05030_),
    .B(_05038_),
    .C(_04891_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10938_ (.A1(_02216_),
    .A2(_02211_),
    .A3(_04949_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10939_ (.A1(_02224_),
    .A2(_05040_),
    .Z(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10940_ (.A1(_04806_),
    .A2(_05041_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10941_ (.A1(_04916_),
    .A2(_05028_),
    .B(_05042_),
    .C(_03816_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10942_ (.A1(_04668_),
    .A2(_05037_),
    .B(_05039_),
    .C(_05043_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10943_ (.A1(_04242_),
    .A2(_04988_),
    .B(_04395_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10944_ (.A1(_04255_),
    .A2(_04270_),
    .A3(_04988_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10945_ (.A1(_04897_),
    .A2(_05046_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10946_ (.A1(_04226_),
    .A2(_05028_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10947_ (.A1(_05045_),
    .A2(_05047_),
    .B(_05048_),
    .C(_04904_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10948_ (.A1(_04333_),
    .A2(_05044_),
    .B(_05049_),
    .C(_00673_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10949_ (.A1(_05035_),
    .A2(_05050_),
    .B(_04948_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10950_ (.A1(_01926_),
    .A2(_04622_),
    .B1(_05033_),
    .B2(_03666_),
    .C(_00882_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10951_ (.A1(_03662_),
    .A2(_05028_),
    .B1(_05051_),
    .B2(_05052_),
    .C(_03832_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10952_ (.A1(\as2650.ivec[7] ),
    .A2(_04972_),
    .B1(_04941_),
    .B2(_05028_),
    .C(_04643_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10953_ (.A1(_05026_),
    .A2(_04700_),
    .B1(_05053_),
    .B2(_05054_),
    .C(_00727_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10954_ (.I(net69),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10955_ (.A1(net69),
    .A2(_05031_),
    .Z(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10956_ (.I(_05056_),
    .Z(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10957_ (.I(_05057_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10958_ (.A1(_04814_),
    .A2(_05046_),
    .B1(_05057_),
    .B2(_04794_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10959_ (.A1(_02229_),
    .A2(_00628_),
    .B(_00779_),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10960_ (.A1(_04811_),
    .A2(_05057_),
    .B(_05060_),
    .C(_00786_),
    .ZN(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10961_ (.A1(_00784_),
    .A2(_00681_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10962_ (.A1(_01155_),
    .A2(_05062_),
    .B(_02331_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10963_ (.A1(_05025_),
    .A2(_05040_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10964_ (.A1(_02229_),
    .A2(_05064_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10965_ (.A1(_02229_),
    .A2(_05064_),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10966_ (.A1(_00444_),
    .A2(_05066_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10967_ (.A1(_04802_),
    .A2(_05056_),
    .B1(_05065_),
    .B2(_05067_),
    .C(_02350_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10968_ (.A1(_05061_),
    .A2(_05063_),
    .B(_05068_),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10969_ (.A1(_05055_),
    .A2(_04228_),
    .B(_02331_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10970_ (.A1(_03749_),
    .A2(_05058_),
    .B(_05070_),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10971_ (.A1(_00783_),
    .A2(_05069_),
    .B1(_05071_),
    .B2(_04364_),
    .C(_04554_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10972_ (.A1(_00522_),
    .A2(_05059_),
    .B(_05072_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10973_ (.A1(_01953_),
    .A2(_04995_),
    .B1(_05057_),
    .B2(_03667_),
    .C(_05073_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10974_ (.A1(_04532_),
    .A2(_05058_),
    .B1(_05074_),
    .B2(_03757_),
    .C(_04744_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10975_ (.I(_04404_),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10976_ (.A1(_05055_),
    .A2(_04701_),
    .B(_05075_),
    .C(_05076_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10977_ (.I(_02235_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10978_ (.A1(_05055_),
    .A2(_05031_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10979_ (.A1(net71),
    .A2(_05078_),
    .Z(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10980_ (.I(_05079_),
    .Z(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10981_ (.A1(_04595_),
    .A2(_05078_),
    .B(_05067_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10982_ (.A1(_02235_),
    .A2(_05081_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10983_ (.A1(_00622_),
    .A2(_00699_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10984_ (.A1(_02235_),
    .A2(_00808_),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10985_ (.A1(_00804_),
    .A2(_05079_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10986_ (.A1(_00805_),
    .A2(_05084_),
    .B(_05085_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10987_ (.A1(_04400_),
    .A2(_05083_),
    .B1(_05086_),
    .B2(_00586_),
    .C(_02901_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10988_ (.A1(_04439_),
    .A2(_05082_),
    .B(_05087_),
    .C(_04904_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10989_ (.A1(_04897_),
    .A2(_05080_),
    .B(_04332_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10990_ (.A1(_04863_),
    .A2(_05089_),
    .B(_03737_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10991_ (.A1(_03816_),
    .A2(_05080_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10992_ (.A1(_04439_),
    .A2(_05084_),
    .B(_05091_),
    .C(_04364_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10993_ (.A1(_05088_),
    .A2(_05090_),
    .B(_03755_),
    .C(_05092_),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10994_ (.A1(_04535_),
    .A2(_05080_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10995_ (.A1(_01974_),
    .A2(_04995_),
    .B(_05093_),
    .C(_05094_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10996_ (.A1(_04532_),
    .A2(_05080_),
    .B1(_05095_),
    .B2(_03757_),
    .C(_04744_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10997_ (.A1(_05077_),
    .A2(_04701_),
    .B(_05096_),
    .C(_05076_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10998_ (.A1(_00799_),
    .A2(_05671_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10999_ (.A1(_02841_),
    .A2(_02772_),
    .B1(_05097_),
    .B2(_00951_),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11000_ (.A1(_01091_),
    .A2(_02723_),
    .B(_00679_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11001_ (.A1(_00451_),
    .A2(_05098_),
    .B1(_05099_),
    .B2(_00866_),
    .C(_00754_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11002_ (.A1(_00725_),
    .A2(_00866_),
    .A3(_03766_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11003_ (.A1(_00864_),
    .A2(_03648_),
    .A3(_03686_),
    .A4(_05101_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11004_ (.A1(_03243_),
    .A2(_00657_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11005_ (.A1(_02607_),
    .A2(_00598_),
    .A3(_05103_),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _11006_ (.A1(_00766_),
    .A2(_00648_),
    .A3(_00870_),
    .A4(_05104_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _11007_ (.A1(_02568_),
    .A2(_02731_),
    .A3(_02739_),
    .A4(_05105_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11008_ (.A1(_05102_),
    .A2(_05106_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11009_ (.A1(_02349_),
    .A2(_00599_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11010_ (.A1(_02746_),
    .A2(_00502_),
    .A3(_03638_),
    .A4(_05108_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11011_ (.A1(_00941_),
    .A2(_02759_),
    .B(_00637_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11012_ (.A1(_00533_),
    .A2(_00973_),
    .A3(_00986_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11013_ (.A1(_00722_),
    .A2(_00979_),
    .B(_05111_),
    .C(_01130_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11014_ (.A1(_03650_),
    .A2(_01131_),
    .A3(_05110_),
    .B1(_05112_),
    .B2(_00555_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11015_ (.A1(_00864_),
    .A2(_05113_),
    .B(_02806_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11016_ (.A1(_00880_),
    .A2(_05109_),
    .B(_05114_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11017_ (.A1(_05100_),
    .A2(_05107_),
    .A3(_05115_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11018_ (.A1(_00963_),
    .A2(_04319_),
    .B(_03745_),
    .C(_00647_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11019_ (.I(_05117_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11020_ (.A1(_03646_),
    .A2(_00904_),
    .B(_02349_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11021_ (.A1(_03646_),
    .A2(_04309_),
    .B1(_05119_),
    .B2(_00959_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11022_ (.A1(_00864_),
    .A2(_04379_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11023_ (.A1(_05120_),
    .A2(_05121_),
    .B(_02742_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11024_ (.A1(_02734_),
    .A2(_05118_),
    .A3(_05122_),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11025_ (.A1(_02763_),
    .A2(_02766_),
    .A3(_05116_),
    .A4(_05123_),
    .Z(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11026_ (.I(_05124_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11027_ (.A1(_03794_),
    .A2(_01012_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11028_ (.A1(_04409_),
    .A2(_01019_),
    .B(_05126_),
    .C(_00971_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11029_ (.A1(_00971_),
    .A2(_01097_),
    .B(_05127_),
    .C(_03781_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11030_ (.I(_05103_),
    .Z(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11031_ (.A1(_00851_),
    .A2(_00872_),
    .A3(_00845_),
    .Z(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11032_ (.I(_05130_),
    .Z(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11033_ (.A1(net78),
    .A2(_05131_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11034_ (.A1(_02028_),
    .A2(_02589_),
    .B(_02724_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11035_ (.I(_05103_),
    .Z(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11036_ (.I(_00847_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11037_ (.A1(_05135_),
    .A2(_04553_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11038_ (.A1(_05132_),
    .A2(_05133_),
    .B(_05134_),
    .C(_05136_),
    .ZN(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11039_ (.I(_00613_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11040_ (.A1(_05129_),
    .A2(_01111_),
    .B(_05137_),
    .C(_05138_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11041_ (.I(_02812_),
    .Z(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11042_ (.A1(_02819_),
    .A2(_01032_),
    .B(_05139_),
    .C(_05140_),
    .ZN(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11043_ (.I(_02764_),
    .Z(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11044_ (.A1(_01277_),
    .A2(_02813_),
    .B(_05141_),
    .C(_05142_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11045_ (.A1(_02845_),
    .A2(_02842_),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11046_ (.A1(_00760_),
    .A2(_05143_),
    .A3(_05144_),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11047_ (.A1(_00428_),
    .A2(_00680_),
    .B1(_02867_),
    .B2(_01139_),
    .C(_00823_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11048_ (.A1(_05128_),
    .A2(_05145_),
    .A3(_05146_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11049_ (.I(_05124_),
    .Z(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11050_ (.A1(_02131_),
    .A2(_01990_),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11051_ (.A1(_01992_),
    .A2(_05149_),
    .Z(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11052_ (.I(_05150_),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11053_ (.I(_05151_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11054_ (.I(_01855_),
    .Z(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11055_ (.I(_01937_),
    .Z(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11056_ (.A1(\as2650.stack[5][0] ),
    .A2(_05153_),
    .B1(_05154_),
    .B2(\as2650.stack[7][0] ),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11057_ (.I(_01940_),
    .Z(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11058_ (.I(_01942_),
    .Z(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11059_ (.A1(_02131_),
    .A2(_01990_),
    .Z(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11060_ (.I(_05158_),
    .Z(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11061_ (.I(_05159_),
    .Z(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11062_ (.A1(\as2650.stack[6][0] ),
    .A2(_05156_),
    .B1(_05157_),
    .B2(\as2650.stack[4][0] ),
    .C(_05160_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11063_ (.I(_01870_),
    .Z(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11064_ (.I(_01941_),
    .Z(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11065_ (.A1(_01771_),
    .A2(_01768_),
    .Z(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11066_ (.I(_05164_),
    .Z(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11067_ (.A1(\as2650.stack[2][0] ),
    .A2(_01940_),
    .B1(_01942_),
    .B2(\as2650.stack[0][0] ),
    .C(_05165_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11068_ (.I(_05166_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11069_ (.A1(\as2650.stack[1][0] ),
    .A2(_05162_),
    .B1(_05163_),
    .B2(\as2650.stack[3][0] ),
    .C(_05167_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11070_ (.A1(_05155_),
    .A2(_05161_),
    .B(_05168_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11071_ (.I(_05151_),
    .Z(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11072_ (.I(_01812_),
    .Z(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11073_ (.I(_01819_),
    .Z(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11074_ (.A1(\as2650.stack[9][0] ),
    .A2(_05171_),
    .B1(_05172_),
    .B2(\as2650.stack[11][0] ),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11075_ (.I(_05164_),
    .Z(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11076_ (.A1(\as2650.stack[10][0] ),
    .A2(_01959_),
    .B1(_01936_),
    .B2(\as2650.stack[8][0] ),
    .C(_05174_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11077_ (.A1(_05173_),
    .A2(_05175_),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11078_ (.I(_05165_),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11079_ (.I(_01877_),
    .Z(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11080_ (.A1(\as2650.stack[13][0] ),
    .A2(_05178_),
    .B1(_01961_),
    .B2(\as2650.stack[12][0] ),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11081_ (.I(_01811_),
    .Z(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11082_ (.A1(\as2650.stack[14][0] ),
    .A2(_05180_),
    .B1(_01962_),
    .B2(\as2650.stack[15][0] ),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11083_ (.A1(_05177_),
    .A2(_05179_),
    .A3(_05181_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11084_ (.A1(_05176_),
    .A2(_05182_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11085_ (.A1(_05170_),
    .A2(_05183_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11086_ (.I(_00755_),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11087_ (.A1(_05152_),
    .A2(_05169_),
    .B(_05184_),
    .C(_05185_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11088_ (.A1(_05147_),
    .A2(_05148_),
    .A3(_05186_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11089_ (.A1(_01102_),
    .A2(_05125_),
    .B(_05187_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11090_ (.A1(_03974_),
    .A2(_05188_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11091_ (.I(_05124_),
    .Z(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11092_ (.A1(_00805_),
    .A2(_00431_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11093_ (.A1(net79),
    .A2(_02589_),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11094_ (.I(_01724_),
    .Z(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11095_ (.A1(_02027_),
    .A2(_00874_),
    .B(_05191_),
    .C(_05192_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11096_ (.A1(_01725_),
    .A2(_04638_),
    .B(_05193_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11097_ (.A1(_05129_),
    .A2(_05194_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11098_ (.A1(_05129_),
    .A2(_01204_),
    .B(_05195_),
    .C(_02819_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11099_ (.A1(_02813_),
    .A2(_05190_),
    .A3(_05196_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11100_ (.A1(_03148_),
    .A2(_02833_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11101_ (.A1(_02811_),
    .A2(_00760_),
    .A3(_05197_),
    .A4(_05198_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11102_ (.I(_00774_),
    .Z(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11103_ (.A1(_04275_),
    .A2(_01127_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11104_ (.I(_00774_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11105_ (.A1(_03948_),
    .A2(_01161_),
    .B(_05202_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11106_ (.A1(_05200_),
    .A2(_01195_),
    .B1(_05201_),
    .B2(_05203_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11107_ (.A1(_02745_),
    .A2(_04651_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11108_ (.A1(_01146_),
    .A2(_00789_),
    .B1(_05205_),
    .B2(_03138_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11109_ (.A1(_04460_),
    .A2(_03679_),
    .B1(_05204_),
    .B2(_03782_),
    .C(_05206_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11110_ (.A1(_05199_),
    .A2(_05207_),
    .B(_00824_),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11111_ (.I(_05165_),
    .Z(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11112_ (.I(_01914_),
    .Z(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11113_ (.A1(\as2650.stack[4][1] ),
    .A2(_05210_),
    .B1(_05154_),
    .B2(\as2650.stack[7][1] ),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11114_ (.I(_01912_),
    .Z(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11115_ (.A1(\as2650.stack[6][1] ),
    .A2(_05212_),
    .B1(_05153_),
    .B2(\as2650.stack[5][1] ),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11116_ (.A1(_05209_),
    .A2(_05211_),
    .A3(_05213_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11117_ (.I(_05158_),
    .Z(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11118_ (.I(_05215_),
    .Z(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11119_ (.A1(\as2650.stack[1][1] ),
    .A2(_05153_),
    .B1(_05154_),
    .B2(\as2650.stack[3][1] ),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11120_ (.A1(\as2650.stack[2][1] ),
    .A2(_05212_),
    .B1(_05157_),
    .B2(\as2650.stack[0][1] ),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11121_ (.A1(_05216_),
    .A2(_05217_),
    .A3(_05218_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11122_ (.A1(_05214_),
    .A2(_05219_),
    .B(_05152_),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11123_ (.I(_00823_),
    .Z(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11124_ (.I(_05151_),
    .Z(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11125_ (.I(_01761_),
    .Z(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11126_ (.A1(\as2650.stack[9][1] ),
    .A2(_02142_),
    .B1(_05223_),
    .B2(\as2650.stack[11][1] ),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11127_ (.I(_01811_),
    .Z(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11128_ (.I(_01816_),
    .Z(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11129_ (.A1(\as2650.stack[10][1] ),
    .A2(_05225_),
    .B1(_05226_),
    .B2(\as2650.stack[8][1] ),
    .C(_05174_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11130_ (.A1(_05224_),
    .A2(_05227_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11131_ (.A1(\as2650.stack[13][1] ),
    .A2(_02142_),
    .B1(_05226_),
    .B2(\as2650.stack[12][1] ),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11132_ (.A1(\as2650.stack[14][1] ),
    .A2(_05225_),
    .B1(_02002_),
    .B2(\as2650.stack[15][1] ),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11133_ (.A1(_05177_),
    .A2(_05229_),
    .A3(_05230_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11134_ (.A1(_05228_),
    .A2(_05231_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11135_ (.A1(_05222_),
    .A2(_05232_),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11136_ (.A1(_05221_),
    .A2(_05233_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11137_ (.A1(_05220_),
    .A2(_05234_),
    .B(_05148_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11138_ (.A1(_03261_),
    .A2(_05189_),
    .B1(_05208_),
    .B2(_05235_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11139_ (.A1(_03974_),
    .A2(_05236_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11140_ (.A1(_04275_),
    .A2(_01261_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11141_ (.I(_00641_),
    .Z(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11142_ (.A1(_05238_),
    .A2(_01286_),
    .B(_00914_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11143_ (.A1(_00775_),
    .A2(_01249_),
    .B1(_05237_),
    .B2(_05239_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11144_ (.I(_00594_),
    .Z(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11145_ (.A1(_02814_),
    .A2(_00842_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11146_ (.I(_05135_),
    .Z(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11147_ (.A1(_05243_),
    .A2(_04696_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11148_ (.I(_05130_),
    .Z(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11149_ (.A1(_02135_),
    .A2(_05245_),
    .B(_05135_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11150_ (.A1(net49),
    .A2(_05245_),
    .B(_05246_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11151_ (.A1(_05242_),
    .A2(_05244_),
    .A3(_05247_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11152_ (.I(_00842_),
    .Z(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11153_ (.I(_01219_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11154_ (.A1(_03138_),
    .A2(_02815_),
    .B1(_05249_),
    .B2(_05250_),
    .C(_05241_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11155_ (.A1(_01269_),
    .A2(_05241_),
    .B1(_05248_),
    .B2(_05251_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11156_ (.A1(_01150_),
    .A2(_02866_),
    .B1(_03653_),
    .B2(_02851_),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11157_ (.A1(_02841_),
    .A2(_03815_),
    .A3(_05252_),
    .B(_05253_),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11158_ (.A1(_00426_),
    .A2(_00680_),
    .B1(_03782_),
    .B2(_05240_),
    .C(_05254_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11159_ (.A1(\as2650.stack[4][2] ),
    .A2(_05210_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11160_ (.I(_01747_),
    .Z(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11161_ (.A1(\as2650.stack[5][2] ),
    .A2(_05257_),
    .B1(_05223_),
    .B2(\as2650.stack[7][2] ),
    .C1(\as2650.stack[6][2] ),
    .C2(_02387_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11162_ (.A1(_05209_),
    .A2(_05256_),
    .A3(_05258_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11163_ (.A1(\as2650.stack[2][2] ),
    .A2(_05212_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11164_ (.A1(\as2650.stack[1][2] ),
    .A2(_05257_),
    .B1(_02271_),
    .B2(\as2650.stack[0][2] ),
    .C1(_05223_),
    .C2(\as2650.stack[3][2] ),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11165_ (.A1(_05216_),
    .A2(_05260_),
    .A3(_05261_),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11166_ (.A1(_05259_),
    .A2(_05262_),
    .B(_05222_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11167_ (.I(_00755_),
    .Z(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11168_ (.I(_05151_),
    .Z(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11169_ (.I(_01782_),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11170_ (.A1(\as2650.stack[13][2] ),
    .A2(_05266_),
    .B1(_02002_),
    .B2(\as2650.stack[15][2] ),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11171_ (.I(_01811_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11172_ (.I(_01900_),
    .Z(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11173_ (.A1(\as2650.stack[14][2] ),
    .A2(_05268_),
    .B1(_05269_),
    .B2(\as2650.stack[12][2] ),
    .C(_05215_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11174_ (.A1(_05267_),
    .A2(_05270_),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11175_ (.A1(\as2650.stack[9][2] ),
    .A2(_05266_),
    .ZN(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11176_ (.A1(\as2650.stack[8][2] ),
    .A2(_01914_),
    .B1(_01937_),
    .B2(\as2650.stack[11][2] ),
    .C1(\as2650.stack[10][2] ),
    .C2(_01933_),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11177_ (.A1(_05160_),
    .A2(_05272_),
    .A3(_05273_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11178_ (.A1(_05271_),
    .A2(_05274_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11179_ (.A1(_05265_),
    .A2(_05275_),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11180_ (.A1(_05264_),
    .A2(_05276_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11181_ (.I(_05124_),
    .Z(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11182_ (.A1(_00757_),
    .A2(_05255_),
    .B1(_05263_),
    .B2(_05277_),
    .C(_05278_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11183_ (.A1(_03267_),
    .A2(_05125_),
    .B(_05279_),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11184_ (.A1(_03974_),
    .A2(_05280_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11185_ (.I(_00696_),
    .Z(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11186_ (.I(_00680_),
    .Z(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11187_ (.A1(_05238_),
    .A2(_03147_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11188_ (.A1(_03761_),
    .A2(_01303_),
    .B(_05202_),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11189_ (.A1(_05200_),
    .A2(_01350_),
    .B1(_05283_),
    .B2(_05284_),
    .C(_03859_),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11190_ (.A1(_01028_),
    .A2(_05245_),
    .ZN(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11191_ (.A1(_02000_),
    .A2(_00874_),
    .B(_05192_),
    .ZN(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11192_ (.A1(_01725_),
    .A2(_04741_),
    .B1(_05286_),
    .B2(_05287_),
    .C(_05242_),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11193_ (.I(_01363_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11194_ (.A1(_03148_),
    .A2(_02815_),
    .B1(_05249_),
    .B2(_05289_),
    .C(_05241_),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11195_ (.A1(_03149_),
    .A2(_02833_),
    .B1(_05288_),
    .B2(_05290_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11196_ (.A1(_01269_),
    .A2(_02866_),
    .B1(_03653_),
    .B2(_02856_),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11197_ (.A1(_02842_),
    .A2(_03815_),
    .A3(_05291_),
    .B(_05292_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11198_ (.A1(_00439_),
    .A2(_05282_),
    .B(_05285_),
    .C(_05293_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11199_ (.A1(\as2650.stack[5][3] ),
    .A2(_05162_),
    .B1(_05163_),
    .B2(\as2650.stack[7][3] ),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11200_ (.I(_01862_),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11201_ (.I(_01869_),
    .Z(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11202_ (.I(_05159_),
    .Z(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11203_ (.A1(\as2650.stack[6][3] ),
    .A2(_05296_),
    .B1(_05297_),
    .B2(\as2650.stack[4][3] ),
    .C(_05298_),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11204_ (.A1(_05295_),
    .A2(_05299_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11205_ (.A1(\as2650.stack[2][3] ),
    .A2(_05296_),
    .B1(_05297_),
    .B2(\as2650.stack[0][3] ),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11206_ (.I(_01870_),
    .Z(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11207_ (.I(_01863_),
    .Z(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11208_ (.A1(\as2650.stack[1][3] ),
    .A2(_05302_),
    .B1(_05303_),
    .B2(\as2650.stack[3][3] ),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11209_ (.A1(_05216_),
    .A2(_05301_),
    .A3(_05304_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11210_ (.A1(_05300_),
    .A2(_05305_),
    .B(_05222_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11211_ (.A1(\as2650.stack[13][3] ),
    .A2(_05266_),
    .B1(_05172_),
    .B2(\as2650.stack[15][3] ),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11212_ (.A1(\as2650.stack[14][3] ),
    .A2(_05268_),
    .B1(_05269_),
    .B2(\as2650.stack[12][3] ),
    .C(_05215_),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11213_ (.A1(_05307_),
    .A2(_05308_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11214_ (.I(_01879_),
    .Z(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11215_ (.A1(\as2650.stack[8][3] ),
    .A2(_05226_),
    .B1(_05310_),
    .B2(\as2650.stack[11][3] ),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11216_ (.A1(\as2650.stack[10][3] ),
    .A2(_05268_),
    .B1(_05178_),
    .B2(\as2650.stack[9][3] ),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11217_ (.A1(_05160_),
    .A2(_05311_),
    .A3(_05312_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11218_ (.A1(_05309_),
    .A2(_05313_),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11219_ (.A1(_05265_),
    .A2(_05314_),
    .ZN(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11220_ (.A1(_05264_),
    .A2(_05315_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11221_ (.A1(_00757_),
    .A2(_05294_),
    .B1(_05306_),
    .B2(_05316_),
    .C(_05278_),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11222_ (.A1(_03273_),
    .A2(_05125_),
    .B(_05317_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11223_ (.A1(_05281_),
    .A2(_05318_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11224_ (.A1(_04275_),
    .A2(_01429_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11225_ (.A1(_03948_),
    .A2(_01445_),
    .B(_05202_),
    .ZN(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11226_ (.A1(_05200_),
    .A2(_01422_),
    .B1(_05319_),
    .B2(_05320_),
    .C(_03859_),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11227_ (.A1(_02927_),
    .A2(_05130_),
    .B(_00847_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11228_ (.A1(_00955_),
    .A2(_05131_),
    .B(_05322_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11229_ (.A1(_02724_),
    .A2(_04786_),
    .B(_05323_),
    .C(_05134_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11230_ (.A1(_05129_),
    .A2(_02223_),
    .B(_05324_),
    .C(_02818_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11231_ (.A1(_01431_),
    .A2(_05138_),
    .B(_05325_),
    .C(_02960_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11232_ (.A1(_01599_),
    .A2(_05140_),
    .B(_05326_),
    .C(_05142_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11233_ (.A1(_03149_),
    .A2(_02867_),
    .B1(_03679_),
    .B2(_02860_),
    .ZN(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11234_ (.A1(_03815_),
    .A2(_05327_),
    .B(_05328_),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11235_ (.A1(_05813_),
    .A2(_05282_),
    .B(_05321_),
    .C(_05329_),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11236_ (.A1(\as2650.stack[1][4] ),
    .A2(_05162_),
    .B1(_05163_),
    .B2(\as2650.stack[3][4] ),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11237_ (.A1(\as2650.stack[2][4] ),
    .A2(_05296_),
    .B1(_05297_),
    .B2(\as2650.stack[0][4] ),
    .C(_05174_),
    .ZN(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11238_ (.A1(_05331_),
    .A2(_05332_),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11239_ (.A1(\as2650.stack[5][4] ),
    .A2(_05302_),
    .B1(_05163_),
    .B2(\as2650.stack[7][4] ),
    .ZN(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11240_ (.A1(\as2650.stack[6][4] ),
    .A2(_02387_),
    .B1(_02271_),
    .B2(\as2650.stack[4][4] ),
    .C(_05298_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11241_ (.A1(_05334_),
    .A2(_05335_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11242_ (.A1(_05333_),
    .A2(_05336_),
    .B(_05265_),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11243_ (.A1(\as2650.stack[13][4] ),
    .A2(_05266_),
    .B1(_05172_),
    .B2(\as2650.stack[15][4] ),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11244_ (.A1(\as2650.stack[14][4] ),
    .A2(_05180_),
    .B1(_05269_),
    .B2(\as2650.stack[12][4] ),
    .C(_05215_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11245_ (.A1(_05338_),
    .A2(_05339_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11246_ (.A1(\as2650.stack[10][4] ),
    .A2(_05225_),
    .B1(_05178_),
    .B2(\as2650.stack[9][4] ),
    .ZN(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11247_ (.A1(\as2650.stack[8][4] ),
    .A2(_01961_),
    .B1(_05310_),
    .B2(\as2650.stack[11][4] ),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11248_ (.A1(_05160_),
    .A2(_05341_),
    .A3(_05342_),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11249_ (.A1(_05340_),
    .A2(_05343_),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11250_ (.A1(_05170_),
    .A2(_05344_),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11251_ (.A1(_05264_),
    .A2(_05345_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11252_ (.A1(_00757_),
    .A2(_05330_),
    .B1(_05337_),
    .B2(_05346_),
    .C(_05278_),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11253_ (.A1(_03279_),
    .A2(_05125_),
    .B(_05347_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11254_ (.A1(_05281_),
    .A2(_05348_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11255_ (.A1(_04129_),
    .A2(_01474_),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11256_ (.A1(_04409_),
    .A2(_01458_),
    .B(_00914_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11257_ (.A1(_00775_),
    .A2(_01501_),
    .B1(_05349_),
    .B2(_05350_),
    .C(_03813_),
    .ZN(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11258_ (.A1(net52),
    .A2(_00873_),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11259_ (.A1(_02610_),
    .A2(_05130_),
    .B(_00847_),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11260_ (.A1(_05352_),
    .A2(_05353_),
    .B(_02814_),
    .C(_00842_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11261_ (.A1(_02724_),
    .A2(_04837_),
    .B(_05354_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11262_ (.A1(_03149_),
    .A2(_02814_),
    .ZN(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11263_ (.A1(_05249_),
    .A2(_01518_),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11264_ (.A1(_05355_),
    .A2(_05356_),
    .A3(_05357_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11265_ (.A1(_02812_),
    .A2(_05358_),
    .ZN(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11266_ (.A1(_02837_),
    .A2(_02960_),
    .B(_05359_),
    .C(_02810_),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11267_ (.A1(_02613_),
    .A2(_05142_),
    .B(_00759_),
    .C(_05360_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11268_ (.A1(_01463_),
    .A2(_00789_),
    .B1(_05205_),
    .B2(_02835_),
    .C(_05361_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11269_ (.A1(_05351_),
    .A2(_05362_),
    .B(_02805_),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11270_ (.I(_05159_),
    .Z(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11271_ (.A1(\as2650.stack[4][5] ),
    .A2(_05210_),
    .B(_05364_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11272_ (.A1(\as2650.stack[5][5] ),
    .A2(_05302_),
    .B1(_05303_),
    .B2(\as2650.stack[7][5] ),
    .C1(\as2650.stack[6][5] ),
    .C2(_05296_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11273_ (.A1(\as2650.stack[2][5] ),
    .A2(_05225_),
    .ZN(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11274_ (.A1(\as2650.stack[1][5] ),
    .A2(_01934_),
    .B1(_01936_),
    .B2(\as2650.stack[0][5] ),
    .C1(_01937_),
    .C2(\as2650.stack[3][5] ),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11275_ (.A1(_05298_),
    .A2(_05367_),
    .A3(_05368_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11276_ (.A1(_05365_),
    .A2(_05366_),
    .B(_05369_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11277_ (.A1(\as2650.stack[13][5] ),
    .A2(_05171_),
    .B1(_05310_),
    .B2(\as2650.stack[15][5] ),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11278_ (.A1(\as2650.stack[14][5] ),
    .A2(_01933_),
    .B1(_01936_),
    .B2(\as2650.stack[12][5] ),
    .C(_05159_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11279_ (.A1(_05371_),
    .A2(_05372_),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11280_ (.A1(\as2650.stack[11][5] ),
    .A2(_02002_),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11281_ (.A1(\as2650.stack[9][5] ),
    .A2(_01934_),
    .B1(_01914_),
    .B2(\as2650.stack[8][5] ),
    .C1(\as2650.stack[10][5] ),
    .C2(_01912_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11282_ (.A1(_05298_),
    .A2(_05374_),
    .A3(_05375_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11283_ (.A1(_05373_),
    .A2(_05376_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11284_ (.A1(_05170_),
    .A2(_05377_),
    .ZN(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11285_ (.A1(_05152_),
    .A2(_05370_),
    .B(_05378_),
    .C(_05185_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11286_ (.A1(_05189_),
    .A2(_05363_),
    .A3(_05379_),
    .ZN(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11287_ (.A1(_03285_),
    .A2(_05189_),
    .B(_05380_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11288_ (.A1(_05281_),
    .A2(_05381_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11289_ (.A1(_05238_),
    .A2(_04081_),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11290_ (.A1(_03761_),
    .A2(_01619_),
    .B(_05202_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11291_ (.A1(_05200_),
    .A2(_01589_),
    .B1(_05382_),
    .B2(_05383_),
    .C(_03859_),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11292_ (.A1(net53),
    .A2(_05131_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11293_ (.A1(net85),
    .A2(_02589_),
    .B(_01724_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11294_ (.A1(_05385_),
    .A2(_05386_),
    .B(_02818_),
    .C(_05134_),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11295_ (.A1(_05243_),
    .A2(_02804_),
    .B(_05387_),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11296_ (.A1(_01599_),
    .A2(_02818_),
    .B1(_05134_),
    .B2(_02234_),
    .C(_02812_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11297_ (.A1(_05388_),
    .A2(_05389_),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11298_ (.A1(_01602_),
    .A2(_02960_),
    .B(_02810_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11299_ (.A1(_02861_),
    .A2(_02810_),
    .B1(_05390_),
    .B2(_05391_),
    .C(_00759_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11300_ (.A1(_02837_),
    .A2(_05205_),
    .B(_05392_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11301_ (.A1(_05801_),
    .A2(_05282_),
    .B(_05384_),
    .C(_05393_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11302_ (.A1(\as2650.stack[6][6] ),
    .A2(_05156_),
    .B1(_05157_),
    .B2(\as2650.stack[4][6] ),
    .ZN(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11303_ (.A1(\as2650.stack[5][6] ),
    .A2(_05302_),
    .B1(_05303_),
    .B2(\as2650.stack[7][6] ),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11304_ (.A1(_05209_),
    .A2(_05395_),
    .A3(_05396_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11305_ (.A1(\as2650.stack[0][6] ),
    .A2(_05297_),
    .B1(_05303_),
    .B2(\as2650.stack[3][6] ),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11306_ (.A1(\as2650.stack[2][6] ),
    .A2(_05156_),
    .B1(_05257_),
    .B2(\as2650.stack[1][6] ),
    .ZN(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11307_ (.A1(_05364_),
    .A2(_05398_),
    .A3(_05399_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11308_ (.A1(_05397_),
    .A2(_05400_),
    .B(_05265_),
    .ZN(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11309_ (.A1(\as2650.stack[9][6] ),
    .A2(_05171_),
    .B1(_05172_),
    .B2(\as2650.stack[11][6] ),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11310_ (.A1(\as2650.stack[10][6] ),
    .A2(_05180_),
    .B1(_05269_),
    .B2(\as2650.stack[8][6] ),
    .C(_05174_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11311_ (.A1(_05402_),
    .A2(_05403_),
    .ZN(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11312_ (.A1(\as2650.stack[14][6] ),
    .A2(_05268_),
    .B1(_01961_),
    .B2(\as2650.stack[12][6] ),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11313_ (.A1(\as2650.stack[13][6] ),
    .A2(_05171_),
    .B1(_05310_),
    .B2(\as2650.stack[15][6] ),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11314_ (.A1(_05177_),
    .A2(_05405_),
    .A3(_05406_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11315_ (.A1(_05404_),
    .A2(_05407_),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11316_ (.A1(_05170_),
    .A2(_05408_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11317_ (.A1(_05185_),
    .A2(_05409_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11318_ (.A1(_00824_),
    .A2(_05394_),
    .B1(_05401_),
    .B2(_05410_),
    .C(_05278_),
    .ZN(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11319_ (.A1(_03609_),
    .A2(_05189_),
    .B(_05411_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11320_ (.A1(_05281_),
    .A2(_05412_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11321_ (.I(_00756_),
    .Z(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11322_ (.A1(_05238_),
    .A2(_01696_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11323_ (.A1(_04409_),
    .A2(_01693_),
    .B(_00914_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11324_ (.A1(_00775_),
    .A2(_01685_),
    .B1(_05414_),
    .B2(_05415_),
    .C(_03813_),
    .ZN(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11325_ (.A1(_05249_),
    .A2(_03465_),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11326_ (.A1(net77),
    .A2(_05245_),
    .ZN(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11327_ (.A1(_02951_),
    .A2(_00874_),
    .B(_05135_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11328_ (.A1(_02592_),
    .A2(_05242_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11329_ (.A1(_05243_),
    .A2(_02924_),
    .B1(_05418_),
    .B2(_05419_),
    .C(_05420_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11330_ (.I(_05421_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11331_ (.A1(_02817_),
    .A2(_02961_),
    .A3(_05417_),
    .A4(_05422_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11332_ (.A1(_05142_),
    .A2(_00759_),
    .A3(_05423_),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11333_ (.A1(_01029_),
    .A2(_02867_),
    .B1(_03679_),
    .B2(_00810_),
    .ZN(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11334_ (.A1(_05424_),
    .A2(_05425_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11335_ (.A1(_05796_),
    .A2(_05282_),
    .B(_05416_),
    .C(_05426_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11336_ (.A1(\as2650.stack[5][7] ),
    .A2(_05153_),
    .B1(_05154_),
    .B2(\as2650.stack[7][7] ),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11337_ (.A1(\as2650.stack[6][7] ),
    .A2(_05212_),
    .B1(_05157_),
    .B2(\as2650.stack[4][7] ),
    .C(_05364_),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11338_ (.A1(_05428_),
    .A2(_05429_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11339_ (.A1(\as2650.stack[0][7] ),
    .A2(_05210_),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11340_ (.A1(\as2650.stack[1][7] ),
    .A2(_05257_),
    .B1(_05223_),
    .B2(\as2650.stack[3][7] ),
    .C1(\as2650.stack[2][7] ),
    .C2(_02387_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11341_ (.A1(_05216_),
    .A2(_05431_),
    .A3(_05432_),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11342_ (.A1(_05430_),
    .A2(_05433_),
    .B(_05152_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11343_ (.A1(\as2650.stack[9][7] ),
    .A2(_02142_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11344_ (.A1(\as2650.stack[8][7] ),
    .A2(_05226_),
    .B1(_01962_),
    .B2(\as2650.stack[11][7] ),
    .C1(\as2650.stack[10][7] ),
    .C2(_05180_),
    .ZN(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11345_ (.A1(_05364_),
    .A2(_05435_),
    .A3(_05436_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11346_ (.A1(\as2650.stack[12][7] ),
    .A2(_02271_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11347_ (.A1(\as2650.stack[13][7] ),
    .A2(_05178_),
    .B1(_01962_),
    .B2(\as2650.stack[15][7] ),
    .C1(\as2650.stack[14][7] ),
    .C2(_01959_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11348_ (.A1(_05209_),
    .A2(_05438_),
    .A3(_05439_),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11349_ (.A1(_05437_),
    .A2(_05440_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11350_ (.A1(_05222_),
    .A2(_05441_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11351_ (.A1(_05221_),
    .A2(_05442_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11352_ (.A1(_05413_),
    .A2(_05427_),
    .B1(_05434_),
    .B2(_05443_),
    .C(_05148_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11353_ (.A1(_02347_),
    .A2(_05148_),
    .Z(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11354_ (.A1(_02625_),
    .A2(_05444_),
    .A3(_05445_),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11355_ (.I(_05446_),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11356_ (.I(\as2650.r123_2[3][0] ),
    .Z(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11357_ (.I(_05447_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11358_ (.I(\as2650.r123_2[3][1] ),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11359_ (.I(_05448_),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11360_ (.I(\as2650.r123_2[3][2] ),
    .Z(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11361_ (.I(_05449_),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11362_ (.I(\as2650.r123_2[3][3] ),
    .Z(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11363_ (.I(_05450_),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11364_ (.I(\as2650.r123_2[3][4] ),
    .Z(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11365_ (.I(_05451_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11366_ (.I(\as2650.r123_2[3][5] ),
    .Z(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11367_ (.I(_05452_),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11368_ (.I(\as2650.r123_2[3][6] ),
    .Z(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11369_ (.I(_05453_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11370_ (.I(\as2650.r123_2[3][7] ),
    .Z(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11371_ (.I(_05454_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11372_ (.A1(_02030_),
    .A2(_02137_),
    .A3(_02664_),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11373_ (.I(_05455_),
    .Z(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11374_ (.I(_05456_),
    .Z(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11375_ (.A1(\as2650.stack[9][8] ),
    .A2(_05456_),
    .ZN(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11376_ (.A1(_02465_),
    .A2(_02138_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11377_ (.I(_05459_),
    .Z(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11378_ (.I(_05460_),
    .Z(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11379_ (.A1(_02663_),
    .A2(_05457_),
    .B(_05458_),
    .C(_05461_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11380_ (.I(_05455_),
    .Z(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11381_ (.A1(\as2650.stack[9][9] ),
    .A2(_05462_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11382_ (.A1(_02672_),
    .A2(_05457_),
    .B(_05461_),
    .C(_05463_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11383_ (.I(_05455_),
    .Z(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11384_ (.A1(\as2650.stack[9][10] ),
    .A2(_05464_),
    .ZN(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11385_ (.A1(_02675_),
    .A2(_05457_),
    .B(_05461_),
    .C(_05465_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11386_ (.A1(\as2650.stack[9][11] ),
    .A2(_05464_),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11387_ (.A1(_02678_),
    .A2(_05457_),
    .B(_05461_),
    .C(_05466_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11388_ (.I(_05456_),
    .Z(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11389_ (.I(_05460_),
    .Z(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11390_ (.A1(\as2650.stack[9][12] ),
    .A2(_05464_),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11391_ (.A1(_02680_),
    .A2(_05467_),
    .B(_05468_),
    .C(_05469_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11392_ (.A1(\as2650.stack[9][13] ),
    .A2(_05464_),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11393_ (.A1(_02684_),
    .A2(_05467_),
    .B(_05468_),
    .C(_05470_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11394_ (.A1(\as2650.stack[9][14] ),
    .A2(_05456_),
    .ZN(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11395_ (.A1(_02686_),
    .A2(_05467_),
    .B(_05468_),
    .C(_05471_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11396_ (.I(_05459_),
    .Z(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11397_ (.I(_05472_),
    .Z(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11398_ (.A1(_02151_),
    .A2(_05467_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11399_ (.A1(_02003_),
    .A2(_02146_),
    .A3(_02438_),
    .ZN(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11400_ (.I(_05475_),
    .Z(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11401_ (.A1(\as2650.stack[9][0] ),
    .A2(_05476_),
    .B(_05468_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11402_ (.A1(_03542_),
    .A2(_05473_),
    .B1(_05474_),
    .B2(_05477_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11403_ (.I(_05475_),
    .Z(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11404_ (.A1(\as2650.stack[9][1] ),
    .A2(_05478_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11405_ (.I(_05455_),
    .Z(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11406_ (.I(_05460_),
    .Z(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11407_ (.A1(_02364_),
    .A2(_05480_),
    .B(_05481_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11408_ (.A1(_03550_),
    .A2(_05473_),
    .B1(_05479_),
    .B2(_05482_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11409_ (.A1(\as2650.stack[9][2] ),
    .A2(_05478_),
    .ZN(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11410_ (.A1(_02074_),
    .A2(_05480_),
    .B(_05481_),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11411_ (.A1(_03555_),
    .A2(_05473_),
    .B1(_05483_),
    .B2(_05484_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11412_ (.A1(\as2650.stack[9][3] ),
    .A2(_05478_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11413_ (.A1(_02087_),
    .A2(_05462_),
    .B(_05481_),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11414_ (.A1(_03558_),
    .A2(_05473_),
    .B1(_05485_),
    .B2(_05486_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11415_ (.I(_05460_),
    .Z(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11416_ (.A1(_03509_),
    .A2(_05480_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11417_ (.A1(\as2650.stack[9][4] ),
    .A2(_05476_),
    .B(_05481_),
    .ZN(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11418_ (.A1(_03561_),
    .A2(_05487_),
    .B1(_05488_),
    .B2(_05489_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11419_ (.A1(\as2650.stack[9][5] ),
    .A2(_05478_),
    .ZN(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11420_ (.A1(_02110_),
    .A2(_05462_),
    .B(_05472_),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11421_ (.A1(_03565_),
    .A2(_05487_),
    .B1(_05490_),
    .B2(_05491_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11422_ (.A1(\as2650.stack[9][6] ),
    .A2(_05476_),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11423_ (.A1(_02119_),
    .A2(_05462_),
    .B(_05472_),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11424_ (.A1(_03568_),
    .A2(_05487_),
    .B1(_05492_),
    .B2(_05493_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11425_ (.A1(_02184_),
    .A2(_05480_),
    .ZN(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11426_ (.A1(\as2650.stack[9][7] ),
    .A2(_05476_),
    .B(_05472_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11427_ (.A1(_03571_),
    .A2(_05487_),
    .B1(_05494_),
    .B2(_05495_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11428_ (.I(_01107_),
    .Z(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11429_ (.A1(_05496_),
    .A2(_03337_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11430_ (.A1(_00514_),
    .A2(_00997_),
    .Z(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11431_ (.I(_05498_),
    .Z(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11432_ (.A1(_01013_),
    .A2(_00934_),
    .A3(_01055_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _11433_ (.A1(_01137_),
    .A2(_00954_),
    .A3(_05500_),
    .A4(_01292_),
    .ZN(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11434_ (.A1(_05697_),
    .A2(_05501_),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11435_ (.A1(_00640_),
    .A2(_01106_),
    .A3(_05502_),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11436_ (.I(_05503_),
    .Z(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11437_ (.A1(_01721_),
    .A2(_05499_),
    .B1(_05504_),
    .B2(\as2650.r123[2][0] ),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11438_ (.A1(_05497_),
    .A2(_05505_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11439_ (.A1(_05496_),
    .A2(_03374_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11440_ (.A1(_01808_),
    .A2(_05499_),
    .B1(_05504_),
    .B2(\as2650.r123[2][1] ),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11441_ (.A1(_05506_),
    .A2(_05507_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11442_ (.A1(_05496_),
    .A2(_03406_),
    .ZN(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11443_ (.A1(_01295_),
    .A2(_05502_),
    .B1(_05504_),
    .B2(\as2650.r123[2][2] ),
    .ZN(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11444_ (.A1(_05508_),
    .A2(_05509_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11445_ (.A1(_05496_),
    .A2(_03431_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11446_ (.A1(_01889_),
    .A2(_05499_),
    .B1(_05504_),
    .B2(\as2650.r123[2][3] ),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11447_ (.A1(_05510_),
    .A2(_05511_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11448_ (.A1(_01223_),
    .A2(_03454_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11449_ (.I(_05503_),
    .Z(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11450_ (.A1(_01449_),
    .A2(_05499_),
    .B1(_05513_),
    .B2(\as2650.r123[2][4] ),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11451_ (.A1(_05512_),
    .A2(_05514_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11452_ (.A1(_01223_),
    .A2(_03473_),
    .ZN(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11453_ (.A1(_01932_),
    .A2(_05498_),
    .B1(_05513_),
    .B2(\as2650.r123[2][5] ),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11454_ (.A1(_05515_),
    .A2(_05516_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11455_ (.A1(_02089_),
    .A2(_00866_),
    .A3(_00657_),
    .A4(_03100_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11456_ (.A1(_01622_),
    .A2(_05498_),
    .B1(_05513_),
    .B2(\as2650.r123[2][6] ),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11457_ (.A1(_05517_),
    .A2(_03484_),
    .B(_05518_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11458_ (.A1(_01707_),
    .A2(_05502_),
    .B1(_05513_),
    .B2(\as2650.r123[2][7] ),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11459_ (.A1(_05517_),
    .A2(_03491_),
    .B(_05519_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11460_ (.I(_02616_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11461_ (.A1(_02901_),
    .A2(_02844_),
    .Z(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11462_ (.I(_00859_),
    .Z(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11463_ (.A1(_01022_),
    .A2(_05672_),
    .A3(_05522_),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11464_ (.A1(_05520_),
    .A2(_04415_),
    .B1(_05521_),
    .B2(_02028_),
    .C(_05523_),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11465_ (.A1(_04620_),
    .A2(_05524_),
    .B(_05221_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11466_ (.A1(_00450_),
    .A2(_02768_),
    .B(_02754_),
    .C(_02740_),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11467_ (.A1(_00702_),
    .A2(_05526_),
    .B(_02581_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11468_ (.A1(_02578_),
    .A2(_04353_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11469_ (.A1(_00884_),
    .A2(_04349_),
    .A3(_05062_),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11470_ (.A1(_04331_),
    .A2(_00950_),
    .A3(_05529_),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11471_ (.A1(_00461_),
    .A2(_00493_),
    .B(_00518_),
    .C(_02010_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11472_ (.A1(_05530_),
    .A2(_05531_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11473_ (.I(_04525_),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11474_ (.A1(_00740_),
    .A2(_02599_),
    .B1(_05533_),
    .B2(_00519_),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11475_ (.A1(_04524_),
    .A2(_05534_),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11476_ (.A1(_00729_),
    .A2(_05532_),
    .B(_05535_),
    .ZN(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11477_ (.A1(_04346_),
    .A2(_05527_),
    .A3(_05528_),
    .A4(_05536_),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11478_ (.A1(_02565_),
    .A2(_04523_),
    .Z(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11479_ (.A1(_02604_),
    .A2(_05537_),
    .A3(_05538_),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11480_ (.I(_05539_),
    .Z(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11481_ (.A1(_03977_),
    .A2(_05525_),
    .B(_05540_),
    .ZN(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11482_ (.A1(_04652_),
    .A2(_05522_),
    .B(_03666_),
    .C(_05524_),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11483_ (.A1(_05264_),
    .A2(_05542_),
    .B(_03780_),
    .ZN(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11484_ (.A1(_02028_),
    .A2(_05543_),
    .Z(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11485_ (.A1(_01772_),
    .A2(_05541_),
    .B1(_05544_),
    .B2(_05540_),
    .C(_00727_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11486_ (.I(\as2650.r123[3][0] ),
    .Z(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11487_ (.I(_05545_),
    .Z(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11488_ (.I(\as2650.r123[3][1] ),
    .Z(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11489_ (.I(_05546_),
    .Z(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11490_ (.I(\as2650.r123[3][2] ),
    .Z(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11491_ (.I(_05547_),
    .Z(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11492_ (.I(\as2650.r123[3][3] ),
    .Z(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11493_ (.I(_05548_),
    .Z(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11494_ (.I(\as2650.r123[3][4] ),
    .Z(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11495_ (.I(_05549_),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11496_ (.I(\as2650.r123[3][5] ),
    .Z(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11497_ (.I(_05550_),
    .Z(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11498_ (.I(\as2650.r123[3][6] ),
    .Z(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11499_ (.I(_05551_),
    .Z(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11500_ (.I(\as2650.r123[3][7] ),
    .Z(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11501_ (.I(_05552_),
    .Z(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11502_ (.I(_05681_),
    .Z(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11503_ (.A1(_02860_),
    .A2(_00751_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11504_ (.A1(_05553_),
    .A2(_04463_),
    .B(_05554_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11505_ (.A1(_04437_),
    .A2(_00751_),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11506_ (.A1(_04948_),
    .A2(_04463_),
    .B(_05555_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11507_ (.A1(_00823_),
    .A2(_04554_),
    .B(_03779_),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11508_ (.A1(_01990_),
    .A2(_01876_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11509_ (.A1(_01992_),
    .A2(_05557_),
    .Z(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11510_ (.A1(_01986_),
    .A2(_05165_),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11511_ (.A1(_05150_),
    .A2(_05559_),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11512_ (.A1(_00826_),
    .A2(_00846_),
    .ZN(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11513_ (.A1(_01306_),
    .A2(_00859_),
    .B(_05192_),
    .C(_02608_),
    .ZN(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11514_ (.A1(_05561_),
    .A2(_05558_),
    .B(_05562_),
    .ZN(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11515_ (.A1(_02856_),
    .A2(_02770_),
    .B(_05563_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11516_ (.A1(_03641_),
    .A2(_05243_),
    .B(_02570_),
    .ZN(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11517_ (.I(_02746_),
    .Z(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11518_ (.A1(_02571_),
    .A2(_05564_),
    .B1(_05565_),
    .B2(_02780_),
    .C(_05566_),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11519_ (.A1(_02777_),
    .A2(_05560_),
    .B(_05567_),
    .ZN(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11520_ (.A1(_05556_),
    .A2(_05558_),
    .B1(_05568_),
    .B2(_03780_),
    .ZN(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11521_ (.A1(_02618_),
    .A2(_05566_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11522_ (.A1(_00730_),
    .A2(_03639_),
    .ZN(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11523_ (.A1(_04437_),
    .A2(_05570_),
    .A3(_05571_),
    .B(_05539_),
    .ZN(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11524_ (.I0(_05569_),
    .I1(_02001_),
    .S(_05572_),
    .Z(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11525_ (.A1(_02625_),
    .A2(_05573_),
    .Z(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11526_ (.I(_05574_),
    .Z(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11527_ (.I(_05570_),
    .Z(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11528_ (.A1(_04462_),
    .A2(_05575_),
    .A3(_05571_),
    .B(_05540_),
    .ZN(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11529_ (.A1(_02648_),
    .A2(_02152_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11530_ (.A1(_05557_),
    .A2(_05577_),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11531_ (.I(_02777_),
    .Z(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11532_ (.A1(_01986_),
    .A2(_05177_),
    .Z(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11533_ (.A1(_01262_),
    .A2(_05522_),
    .B(_05192_),
    .C(_02350_),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11534_ (.A1(_05561_),
    .A2(_05578_),
    .B(_05581_),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11535_ (.A1(_04462_),
    .A2(_02770_),
    .B(_05582_),
    .ZN(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11536_ (.A1(_04626_),
    .A2(_05565_),
    .B1(_05583_),
    .B2(_02621_),
    .C(_05566_),
    .ZN(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11537_ (.A1(_05579_),
    .A2(_05580_),
    .B(_05584_),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11538_ (.A1(_05556_),
    .A2(_05578_),
    .B1(_05585_),
    .B2(_04298_),
    .ZN(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11539_ (.A1(_05576_),
    .A2(_05586_),
    .B(_04501_),
    .ZN(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11540_ (.A1(_02648_),
    .A2(_05576_),
    .B(_05587_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11541_ (.A1(_04460_),
    .A2(_05575_),
    .A3(_05571_),
    .B(_05540_),
    .ZN(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11542_ (.A1(_01773_),
    .A2(_02153_),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11543_ (.A1(_05156_),
    .A2(_05162_),
    .ZN(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11544_ (.A1(_05672_),
    .A2(_00861_),
    .A3(_05589_),
    .B1(_04429_),
    .B2(_05522_),
    .ZN(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11545_ (.A1(_02847_),
    .A2(_02770_),
    .B(_05591_),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11546_ (.A1(_05590_),
    .A2(_05565_),
    .B1(_05592_),
    .B2(_02621_),
    .C(_05566_),
    .ZN(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11547_ (.A1(_02027_),
    .A2(_05579_),
    .B(_05593_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11548_ (.A1(_05589_),
    .A2(_05556_),
    .B1(_05594_),
    .B2(_04298_),
    .ZN(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11549_ (.A1(_05588_),
    .A2(_05595_),
    .B(_04501_),
    .ZN(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11550_ (.A1(_02027_),
    .A2(_05588_),
    .B(_05596_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11551_ (.A1(_03657_),
    .A2(_05140_),
    .A3(_02768_),
    .B(_01038_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11552_ (.A1(_03657_),
    .A2(_01498_),
    .A3(_02748_),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11553_ (.A1(_05108_),
    .A2(_05598_),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11554_ (.A1(_02756_),
    .A2(_02731_),
    .Z(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11555_ (.A1(_00773_),
    .A2(_01090_),
    .B(_04225_),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _11556_ (.A1(_00736_),
    .A2(_02841_),
    .A3(_00950_),
    .A4(_02735_),
    .ZN(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11557_ (.A1(_00754_),
    .A2(_04621_),
    .B1(_05601_),
    .B2(_02740_),
    .C(_05602_),
    .ZN(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11558_ (.A1(_05600_),
    .A2(_05603_),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _11559_ (.A1(_02584_),
    .A2(_02725_),
    .A3(_02728_),
    .A4(_02774_),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11560_ (.A1(_05599_),
    .A2(_05604_),
    .A3(_05605_),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11561_ (.A1(_00863_),
    .A2(_02732_),
    .A3(_00613_),
    .A4(_05131_),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11562_ (.A1(_00850_),
    .A2(_02768_),
    .B(_02752_),
    .C(_05607_),
    .ZN(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _11563_ (.A1(_00471_),
    .A2(_02757_),
    .A3(_02734_),
    .A4(_05608_),
    .Z(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11564_ (.A1(_02076_),
    .A2(_05597_),
    .B(_05606_),
    .C(_05609_),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11565_ (.A1(_02965_),
    .A2(_05521_),
    .B(_05610_),
    .ZN(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11566_ (.A1(_01576_),
    .A2(_01583_),
    .B(_02875_),
    .C(_01679_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11567_ (.A1(_01327_),
    .A2(_02880_),
    .ZN(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11568_ (.A1(_01674_),
    .A2(_01672_),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11569_ (.A1(_01675_),
    .A2(_05614_),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11570_ (.A1(_05612_),
    .A2(_05613_),
    .B1(_05615_),
    .B2(_00839_),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11571_ (.A1(_02956_),
    .A2(_04416_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11572_ (.A1(_05138_),
    .A2(_04417_),
    .A3(_05617_),
    .ZN(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11573_ (.A1(_02834_),
    .A2(_02819_),
    .B(_05618_),
    .C(_05140_),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11574_ (.A1(_00427_),
    .A2(_02813_),
    .B(_05619_),
    .C(_03661_),
    .ZN(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11575_ (.A1(_04161_),
    .A2(_05616_),
    .B(_05620_),
    .ZN(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11576_ (.A1(_04545_),
    .A2(_04552_),
    .B(_05579_),
    .ZN(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11577_ (.A1(_02778_),
    .A2(_05621_),
    .B(_05611_),
    .C(_05622_),
    .ZN(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11578_ (.A1(_01983_),
    .A2(_05611_),
    .B(_05623_),
    .C(_05076_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11579_ (.A1(_04652_),
    .A2(_02614_),
    .A3(_02965_),
    .B(_05610_),
    .ZN(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _11580_ (.A1(_01327_),
    .A2(_01416_),
    .A3(_01421_),
    .ZN(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11581_ (.A1(_02956_),
    .A2(_02609_),
    .ZN(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11582_ (.A1(_05138_),
    .A2(_04446_),
    .A3(_05626_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11583_ (.A1(_05356_),
    .A2(_05627_),
    .B(_05241_),
    .ZN(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11584_ (.A1(_01462_),
    .A2(_02833_),
    .B(_05628_),
    .C(_04062_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11585_ (.A1(_05553_),
    .A2(_05625_),
    .B(_05629_),
    .C(_00756_),
    .ZN(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11586_ (.A1(_05413_),
    .A2(_04837_),
    .B(_05624_),
    .C(_05630_),
    .ZN(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11587_ (.A1(_02101_),
    .A2(_05624_),
    .B(_05631_),
    .C(_05076_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11588_ (.A1(_03642_),
    .A2(_04462_),
    .A3(_02965_),
    .ZN(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11589_ (.A1(_02746_),
    .A2(_00951_),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11590_ (.A1(_00662_),
    .A2(_05633_),
    .ZN(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _11591_ (.A1(_05608_),
    .A2(_05606_),
    .A3(_05632_),
    .A4(_05634_),
    .ZN(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11592_ (.A1(net49),
    .A2(_05635_),
    .Z(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11593_ (.I0(_01675_),
    .I1(_01674_),
    .S(_01685_),
    .Z(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11594_ (.I(_02956_),
    .Z(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11595_ (.A1(_05638_),
    .A2(_04433_),
    .B(_04435_),
    .C(_05553_),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11596_ (.A1(_05553_),
    .A2(_05637_),
    .B(_05639_),
    .ZN(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11597_ (.A1(_05221_),
    .A2(_04696_),
    .ZN(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11598_ (.A1(_05413_),
    .A2(_05640_),
    .B(_05635_),
    .C(_05641_),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11599_ (.A1(_03972_),
    .A2(_05636_),
    .A3(_05642_),
    .Z(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11600_ (.I(_05643_),
    .Z(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11601_ (.I(_05608_),
    .ZN(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11602_ (.A1(_02764_),
    .A2(_02740_),
    .A3(_03638_),
    .A4(_05633_),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _11603_ (.A1(_02737_),
    .A2(_02569_),
    .A3(_05600_),
    .A4(_05645_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11604_ (.A1(_05599_),
    .A2(_05605_),
    .A3(_05644_),
    .A4(_05646_),
    .Z(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11605_ (.A1(_00824_),
    .A2(_02903_),
    .A3(_02860_),
    .B(_05647_),
    .ZN(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11606_ (.A1(_05638_),
    .A2(_04443_),
    .ZN(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11607_ (.A1(_05579_),
    .A2(_04444_),
    .A3(_05649_),
    .ZN(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11608_ (.A1(_02778_),
    .A2(_04786_),
    .B(_05650_),
    .ZN(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11609_ (.A1(_01290_),
    .A2(_05648_),
    .B1(_05651_),
    .B2(_05647_),
    .ZN(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11610_ (.A1(_00697_),
    .A2(_05652_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11611_ (.A1(_04437_),
    .A2(_05575_),
    .B(_05647_),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11612_ (.A1(_02805_),
    .A2(_04741_),
    .ZN(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11613_ (.A1(_05638_),
    .A2(_04440_),
    .B(_04441_),
    .C(_05185_),
    .ZN(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11614_ (.A1(_05653_),
    .A2(_05654_),
    .A3(_05655_),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11615_ (.A1(_02077_),
    .A2(_05653_),
    .B(_05656_),
    .C(_00712_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11616_ (.A1(_04460_),
    .A2(_05575_),
    .B(_05647_),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11617_ (.A1(_05638_),
    .A2(_04429_),
    .B(_04430_),
    .C(_00756_),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11618_ (.A1(_05413_),
    .A2(_04638_),
    .B(_05657_),
    .C(_05658_),
    .ZN(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11619_ (.A1(_02050_),
    .A2(_05657_),
    .B(_05659_),
    .C(_00712_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11620_ (.A1(_04652_),
    .A2(_04399_),
    .ZN(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11621_ (.A1(_02340_),
    .A2(_05660_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11622_ (.A1(net85),
    .A2(_05661_),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11623_ (.A1(_02616_),
    .A2(_04448_),
    .B(_04449_),
    .C(_05661_),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11624_ (.A1(_03972_),
    .A2(_05663_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11625_ (.A1(_05662_),
    .A2(_05664_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11626_ (.A1(_05674_),
    .A2(_04394_),
    .B(_02340_),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11627_ (.A1(_02616_),
    .A2(_04443_),
    .ZN(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11628_ (.A1(_04444_),
    .A2(_05666_),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11629_ (.A1(net74),
    .A2(_05665_),
    .ZN(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11630_ (.A1(_05665_),
    .A2(_05667_),
    .B(_05668_),
    .C(_00712_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11631_ (.D(_00014_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11632_ (.D(_00015_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11633_ (.D(_00016_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11634_ (.D(_00017_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11635_ (.D(_00018_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11636_ (.D(_00019_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11637_ (.D(_00020_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11638_ (.D(_00021_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11639_ (.D(_00022_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11640_ (.D(_00023_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11641_ (.D(_00024_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11642_ (.D(_00025_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11643_ (.D(_00026_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11644_ (.D(_00027_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11645_ (.D(_00028_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11646_ (.D(_00029_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11647_ (.D(_00030_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11648_ (.D(_00031_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11649_ (.D(_00032_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11650_ (.D(_00033_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11651_ (.D(_00034_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11652_ (.D(_00035_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11653_ (.D(_00036_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11654_ (.D(_00037_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11655_ (.D(_00038_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11656_ (.D(_00039_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11657_ (.D(_00040_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11658_ (.D(_00041_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11659_ (.D(_00042_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11660_ (.D(_00043_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11661_ (.D(_00044_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11662_ (.D(_00045_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11663_ (.D(_00046_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11664_ (.D(_00047_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11665_ (.D(_00048_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11666_ (.D(_00049_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11667_ (.D(_00050_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11668_ (.D(_00051_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11669_ (.D(_00052_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11670_ (.D(_00053_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11671_ (.D(_00054_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11672_ (.D(_00055_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11673_ (.D(_00056_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11674_ (.D(_00057_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11675_ (.D(_00058_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11676_ (.D(_00059_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11677_ (.D(_00060_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11678_ (.D(_00061_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11679_ (.D(_00062_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11680_ (.D(_00063_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11681_ (.D(_00064_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11682_ (.D(_00065_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11683_ (.D(_00066_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11684_ (.D(_00067_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11685_ (.D(_00068_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11686_ (.D(_00069_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11687_ (.D(_00070_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11688_ (.D(_00071_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11689_ (.D(_00072_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11690_ (.D(_00073_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11691_ (.D(_00074_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11692_ (.D(_00075_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11693_ (.D(_00076_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11694_ (.D(_00077_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11695_ (.D(_00078_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11696_ (.D(_00079_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11697_ (.D(_00080_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11698_ (.D(_00081_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11699_ (.D(_00082_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11700_ (.D(_00083_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11701_ (.D(_00084_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11702_ (.D(_00085_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11703_ (.D(_00086_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11704_ (.D(_00087_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11705_ (.D(_00088_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11706_ (.D(_00089_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(net77));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11707_ (.D(_00090_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11708_ (.D(_00091_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11709_ (.D(_00092_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11710_ (.D(_00093_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11711_ (.D(_00094_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11712_ (.D(_00095_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11713_ (.D(_00096_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11714_ (.D(_00097_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11715_ (.D(_00098_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11716_ (.D(_00099_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11717_ (.D(_00100_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11718_ (.D(_00101_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11719_ (.D(_00102_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11720_ (.D(_00103_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11721_ (.D(_00104_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11722_ (.D(_00105_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11723_ (.D(_00106_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11724_ (.D(_00107_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11725_ (.D(_00108_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11726_ (.D(_00109_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11727_ (.D(_00110_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11728_ (.D(_00111_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11729_ (.D(_00112_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11730_ (.D(_00113_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11731_ (.D(_00114_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11732_ (.D(_00115_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11733_ (.D(_00116_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11734_ (.D(_00117_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11735_ (.D(_00118_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11736_ (.D(_00119_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11737_ (.D(_00120_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11738_ (.D(_00121_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11739_ (.D(_00122_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11740_ (.D(_00123_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11741_ (.D(_00124_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11742_ (.D(_00125_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11743_ (.D(_00126_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11744_ (.D(_00127_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11745_ (.D(_00128_),
    .CLK(clknet_4_8_0_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11746_ (.D(_00129_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11747_ (.D(_00130_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11748_ (.D(_00131_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11749_ (.D(_00132_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11750_ (.D(_00133_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11751_ (.D(_00134_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11752_ (.D(_00135_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11753_ (.D(_00136_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11754_ (.D(_00137_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11755_ (.D(_00138_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11756_ (.D(_00139_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11757_ (.D(_00140_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11758_ (.D(_00141_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11759_ (.D(_00142_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11760_ (.D(_00143_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11761_ (.D(_00144_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11762_ (.D(_00145_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11763_ (.D(_00146_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11764_ (.D(_00147_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11765_ (.D(_00148_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11766_ (.D(_00149_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net75));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11767_ (.D(_00150_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11768_ (.D(_00151_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11769_ (.D(_00152_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11770_ (.D(_00153_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11771_ (.D(_00154_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11772_ (.D(_00155_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11773_ (.D(_00156_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11774_ (.D(_00157_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11775_ (.D(_00158_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11776_ (.D(_00159_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11777_ (.D(_00160_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11778_ (.D(_00161_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11779_ (.D(_00162_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11780_ (.D(_00163_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11781_ (.D(_00164_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11782_ (.D(_00165_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11783_ (.D(_00166_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11784_ (.D(_00167_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11785_ (.D(_00168_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11786_ (.D(_00169_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11787_ (.D(_00170_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11788_ (.D(_00171_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11789_ (.D(_00172_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11790_ (.D(_00173_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11791_ (.D(_00174_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11792_ (.D(_00175_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11793_ (.D(_00176_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11794_ (.D(_00177_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11795_ (.D(_00178_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11796_ (.D(_00179_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11797_ (.D(_00180_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11798_ (.D(_00181_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11799_ (.D(_00182_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11800_ (.D(_00183_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11801_ (.D(_00184_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11802_ (.D(_00185_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net53));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11803_ (.D(_00186_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net54));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11804_ (.D(_00187_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11805_ (.D(_00188_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11806_ (.D(_00189_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11807_ (.D(_00190_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11808_ (.D(_00191_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11809_ (.D(_00192_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11810_ (.D(_00193_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11811_ (.D(_00194_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11812_ (.D(_00195_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11813_ (.D(_00196_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11814_ (.D(_00197_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11815_ (.D(_00198_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11816_ (.D(_00199_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11817_ (.D(_00200_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11818_ (.D(_00201_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11819_ (.D(_00202_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11820_ (.D(_00203_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11821_ (.D(_00204_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11822_ (.D(_00205_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11823_ (.D(_00206_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11824_ (.D(_00207_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11825_ (.D(_00208_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11826_ (.D(_00209_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11827_ (.D(_00210_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11828_ (.D(_00211_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11829_ (.D(_00212_),
    .CLK(clknet_4_7_0_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11830_ (.D(_00213_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11831_ (.D(_00214_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11832_ (.D(_00215_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11833_ (.D(_00216_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11834_ (.D(_00217_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11835_ (.D(_00218_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11836_ (.D(_00219_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11837_ (.D(_00220_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11838_ (.D(_00221_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11839_ (.D(_00222_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11840_ (.D(_00223_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11841_ (.D(_00224_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11842_ (.D(_00225_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11843_ (.D(_00226_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11844_ (.D(_00000_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11845_ (.D(_00005_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11846_ (.D(_00006_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11847_ (.D(_00007_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11848_ (.D(_00008_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11849_ (.D(_00009_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11850_ (.D(_00010_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11851_ (.D(_00011_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11852_ (.D(_00012_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11853_ (.D(_00013_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11854_ (.D(_00001_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11855_ (.D(_00002_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11856_ (.D(_00003_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.cycle[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11857_ (.D(_00004_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\as2650.cycle[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11858_ (.D(_00227_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11859_ (.D(_00228_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11860_ (.D(_00229_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11861_ (.D(_00230_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11862_ (.D(_00231_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11863_ (.D(_00232_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11864_ (.D(_00233_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11865_ (.D(_00234_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11866_ (.D(_00235_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11867_ (.D(_00236_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11868_ (.D(_00237_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11869_ (.D(_00238_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11870_ (.D(_00239_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11871_ (.D(_00240_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11872_ (.D(_00241_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11873_ (.D(_00242_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11874_ (.D(_00243_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11875_ (.D(_00244_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11876_ (.D(_00245_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11877_ (.D(_00246_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11878_ (.D(_00247_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11879_ (.D(_00248_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11880_ (.D(_00249_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11881_ (.D(_00250_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11882_ (.D(_00251_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11883_ (.D(_00252_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11884_ (.D(_00253_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11885_ (.D(_00254_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11886_ (.D(_00255_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11887_ (.D(_00256_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11888_ (.D(_00257_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11889_ (.D(_00258_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11890_ (.D(_00259_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11891_ (.D(_00260_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11892_ (.D(_00261_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11893_ (.D(_00262_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11894_ (.D(_00263_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11895_ (.D(_00264_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11896_ (.D(_00265_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11897_ (.D(_00266_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11898_ (.D(_00267_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11899_ (.D(_00268_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11900_ (.D(_00269_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11901_ (.D(_00270_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11902_ (.D(_00271_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11903_ (.D(_00272_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11904_ (.D(_00273_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11905_ (.D(_00274_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11906_ (.D(_00275_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.ivec[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11907_ (.D(_00276_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.ivec[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11908_ (.D(_00277_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.ivec[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11909_ (.D(_00278_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.ivec[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11910_ (.D(_00279_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.ivec[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11911_ (.D(_00280_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.ivec[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11912_ (.D(_00281_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.ivec[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11913_ (.D(_00282_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.ivec[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11914_ (.D(_00283_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11915_ (.D(_00284_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11916_ (.D(_00285_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11917_ (.D(_00286_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11918_ (.D(_00287_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11919_ (.D(_00288_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11920_ (.D(_00289_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11921_ (.D(_00290_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11922_ (.D(_00291_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11923_ (.D(_00292_),
    .CLK(clknet_4_6_0_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11924_ (.D(_00293_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11925_ (.D(_00294_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11926_ (.D(_00295_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11927_ (.D(_00296_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11928_ (.D(_00297_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11929_ (.D(_00298_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11930_ (.D(_00299_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11931_ (.D(_00300_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11932_ (.D(_00301_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11933_ (.D(_00302_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11934_ (.D(_00303_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11935_ (.D(_00304_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11936_ (.D(_00305_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11937_ (.D(_00306_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11938_ (.D(_00307_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11939_ (.D(_00308_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11940_ (.D(_00309_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11941_ (.D(_00310_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11942_ (.D(_00311_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11943_ (.D(_00312_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11944_ (.D(_00313_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11945_ (.D(_00314_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11946_ (.D(_00315_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11947_ (.D(_00316_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11948_ (.D(_00317_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(\as2650.last_intr ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11949_ (.D(_00318_),
    .CLK(clknet_4_6_0_wb_clk_i),
    .Q(\as2650.prefixed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11950_ (.D(_00319_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11951_ (.D(_00320_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11952_ (.D(_00321_),
    .CLK(clknet_4_5_0_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11953_ (.D(_00322_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11954_ (.D(_00323_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11955_ (.D(_00324_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11956_ (.D(_00325_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11957_ (.D(_00326_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11958_ (.D(_00327_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11959_ (.D(_00328_),
    .CLK(clknet_4_5_0_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11960_ (.D(_00329_),
    .CLK(clknet_4_7_0_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11961_ (.D(_00330_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11962_ (.D(_00331_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11963_ (.D(_00332_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11964_ (.D(_00333_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.alu_op[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11965_ (.D(_00334_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11966_ (.D(_00335_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net72));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11967_ (.D(_00336_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11968_ (.D(_00337_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11969_ (.D(_00338_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11970_ (.D(_00339_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net46));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11971_ (.D(_00340_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net47));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11972_ (.D(_00341_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11973_ (.D(_00342_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11974_ (.D(_00343_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11975_ (.D(_00344_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(net55));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11976_ (.D(_00345_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(net56));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11977_ (.D(_00346_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(net57));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11978_ (.D(_00347_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(net58));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11979_ (.D(_00348_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(net60));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11980_ (.D(_00349_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(net61));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11981_ (.D(_00350_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(net62));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11982_ (.D(_00351_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(net63));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11983_ (.D(_00352_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net64));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11984_ (.D(_00353_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net65));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11985_ (.D(_00354_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11986_ (.D(_00355_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11987_ (.D(_00356_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net68));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11988_ (.D(_00357_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(net69));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11989_ (.D(_00358_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(net71));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11990_ (.D(_00359_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11991_ (.D(_00360_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11992_ (.D(_00361_),
    .CLK(clknet_4_5_0_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11993_ (.D(_00362_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11994_ (.D(_00363_),
    .CLK(clknet_4_5_0_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11995_ (.D(_00364_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11996_ (.D(_00365_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11997_ (.D(_00366_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11998_ (.D(_00367_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.r123_2[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11999_ (.D(_00368_),
    .CLK(clknet_4_15_0_wb_clk_i),
    .Q(\as2650.r123_2[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12000_ (.D(_00369_),
    .CLK(clknet_4_10_0_wb_clk_i),
    .Q(\as2650.r123_2[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12001_ (.D(_00370_),
    .CLK(clknet_opt_2_0_wb_clk_i),
    .Q(\as2650.r123_2[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12002_ (.D(_00371_),
    .CLK(clknet_4_15_0_wb_clk_i),
    .Q(\as2650.r123_2[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12003_ (.D(_00372_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123_2[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12004_ (.D(_00373_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.r123_2[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12005_ (.D(_00374_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.r123_2[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12006_ (.D(_00375_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12007_ (.D(_00376_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(\as2650.stack[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12008_ (.D(_00377_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12009_ (.D(_00378_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12010_ (.D(_00379_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12011_ (.D(_00380_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12012_ (.D(_00381_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(\as2650.stack[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12013_ (.D(_00382_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12014_ (.D(_00383_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12015_ (.D(_00384_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12016_ (.D(_00385_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12017_ (.D(_00386_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12018_ (.D(_00387_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12019_ (.D(_00388_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12020_ (.D(_00389_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12021_ (.D(_00390_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12022_ (.D(_00391_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12023_ (.D(_00392_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12024_ (.D(_00393_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12025_ (.D(_00394_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12026_ (.D(_00395_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12027_ (.D(_00396_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12028_ (.D(_00397_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12029_ (.D(_00398_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(net48));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12030_ (.D(_00399_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12031_ (.D(_00400_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12032_ (.D(_00401_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12033_ (.D(_00402_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12034_ (.D(_00403_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12035_ (.D(_00404_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12036_ (.D(_00405_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12037_ (.D(_00406_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12038_ (.D(_00407_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12039_ (.D(_00408_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12040_ (.D(_00409_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(net73));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12041_ (.D(_00410_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(net70));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12042_ (.D(_00411_),
    .CLK(clknet_opt_1_0_wb_clk_i),
    .Q(net59));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12043_ (.D(_00412_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(net78));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12044_ (.D(_00413_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(net52));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12045_ (.D(_00414_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(net49));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12046_ (.D(_00415_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net51));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12047_ (.D(_00416_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(net50));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12048_ (.D(_00417_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(net79));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12049_ (.D(_00418_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12050_ (.D(_00419_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(net74));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_142 (.Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_143 (.Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_144 (.Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_145 (.Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_146 (.Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_147 (.Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_148 (.Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_149 (.Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_150 (.Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_151 (.Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_152 (.Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_153 (.Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_154 (.Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_155 (.Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_156 (.Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_157 (.Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_158 (.Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_159 (.Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_160 (.Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_161 (.Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_162 (.Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_163 (.Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_164 (.Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_165 (.Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_166 (.Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_167 (.Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_141 (.Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12124_ (.I(net80),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12125_ (.I(net80),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12126_ (.I(net80),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12127_ (.I(net80),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12128_ (.I(net81),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12129_ (.I(net81),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12130_ (.I(net81),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12131_ (.I(net85),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(io_in[33]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(io_in[34]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(io_in[35]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(io_in[5]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input9 (.I(io_in[6]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(io_in[7]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(io_in[8]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input12 (.I(io_in[9]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net13),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net84),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output46 (.I(net46),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output47 (.I(net47),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output48 (.I(net48),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output49 (.I(net49),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output50 (.I(net50),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output51 (.I(net51),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output52 (.I(net52),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output53 (.I(net94),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output54 (.I(net54),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output55 (.I(net90),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output56 (.I(net56),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output57 (.I(net89),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output58 (.I(net58),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output59 (.I(net86),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output60 (.I(net60),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output61 (.I(net61),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output62 (.I(net62),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output63 (.I(net63),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output64 (.I(net88),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output65 (.I(net87),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output66 (.I(net66),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output67 (.I(net67),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output68 (.I(net68),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output69 (.I(net69),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output70 (.I(net70),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output71 (.I(net71),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output72 (.I(net72),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output73 (.I(net73),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output74 (.I(net74),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output75 (.I(net75),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output76 (.I(net76),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output77 (.I(net77),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output78 (.I(net78),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output79 (.I(net79),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout80 (.I(net82),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout81 (.I(net82),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout82 (.I(net83),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout83 (.I(net84),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout84 (.I(net15),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout85 (.I(net29),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout86 (.I(net59),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout87 (.I(net65),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout88 (.I(net64),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout89 (.I(net57),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout90 (.I(net55),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout91 (.I(net27),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout92 (.I(net42),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout93 (.I(net30),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout94 (.I(net53),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_4_14_0_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_4_14_0_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_4_14_0_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_84_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_90_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_91_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_93_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_95_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_98_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_104_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_107_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_109_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_112_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_119_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_125_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_126_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_127_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_128_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_129_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_130_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_131_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_131_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_132_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_133_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_135_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_15_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_0_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11855__D (.I(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11845__D (.I(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11847__D (.I(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__D (.I(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11850__D (.I(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11636__D (.I(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__D (.I(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__D (.I(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11706__D (.I(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__D (.I(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11721__D (.I(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__D (.I(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11809__D (.I(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11818__D (.I(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11825__D (.I(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__D (.I(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11922__D (.I(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11925__D (.I(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11926__D (.I(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11927__D (.I(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11928__D (.I(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11929__D (.I(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11930__D (.I(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11931__D (.I(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11932__D (.I(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11938__D (.I(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11960__D (.I(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11961__D (.I(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11990__D (.I(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11991__D (.I(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11992__D (.I(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11994__D (.I(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11995__D (.I(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11996__D (.I(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12029__D (.I(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__D (.I(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12041__D (.I(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A1 (.I(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05963__A2 (.I(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__A1 (.I(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__A1 (.I(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__I (.I(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__A1 (.I(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A1 (.I(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__A1 (.I(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__A1 (.I(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__A2 (.I(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__A1 (.I(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A2 (.I(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__A1 (.I(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__A2 (.I(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A1 (.I(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__A1 (.I(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__A1 (.I(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A3 (.I(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__A2 (.I(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__A3 (.I(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__A2 (.I(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A2 (.I(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A2 (.I(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__I (.I(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__B (.I(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A3 (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__I1 (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A1 (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__A2 (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__A1 (.I(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__A1 (.I(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__I (.I(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05980__A1 (.I(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A1 (.I(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A1 (.I(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__A1 (.I(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__A4 (.I(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__S (.I(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__A3 (.I(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A1 (.I(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05984__A2 (.I(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__I (.I(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__I (.I(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A1 (.I(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__I (.I(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10693__I (.I(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05986__I (.I(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__A1 (.I(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A1 (.I(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__B2 (.I(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__A2 (.I(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__A2 (.I(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A2 (.I(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__I (.I(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__I (.I(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__I (.I(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A1 (.I(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__A2 (.I(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__A1 (.I(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__A2 (.I(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__A1 (.I(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__I (.I(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__A1 (.I(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__A2 (.I(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__A2 (.I(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__I (.I(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__A1 (.I(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__I (.I(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__I (.I(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__I (.I(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10831__A1 (.I(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__B2 (.I(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__A1 (.I(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__A3 (.I(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__A2 (.I(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06056__I (.I(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__A2 (.I(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A2 (.I(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__A2 (.I(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__I (.I(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A2 (.I(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__I (.I(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A1 (.I(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__A1 (.I(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A1 (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A1 (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__I (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__A1 (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A1 (.I(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__A1 (.I(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__A1 (.I(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__A1 (.I(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__A1 (.I(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A2 (.I(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06514__A2 (.I(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__A2 (.I(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__A1 (.I(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A2 (.I(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__A2 (.I(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A4 (.I(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A2 (.I(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__A1 (.I(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__A3 (.I(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A1 (.I(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A1 (.I(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__A2 (.I(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__I (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__I (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__A1 (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__A1 (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__B (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A1 (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__A1 (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06010__A1 (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__A1 (.I(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__A1 (.I(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__A1 (.I(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06010__A2 (.I(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A2 (.I(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A1 (.I(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__I (.I(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A1 (.I(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07589__A1 (.I(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__I (.I(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__A2 (.I(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11563__A1 (.I(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A1 (.I(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__A2 (.I(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A1 (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__A1 (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A1 (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__A2 (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__B2 (.I(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__I (.I(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__I (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__A1 (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06392__A1 (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__A1 (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__A1 (.I(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__I (.I(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__A2 (.I(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A1 (.I(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__I (.I(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__A1 (.I(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__I (.I(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__A1 (.I(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A1 (.I(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A2 (.I(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__A2 (.I(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__A1 (.I(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__A2 (.I(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A1 (.I(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__A1 (.I(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A2 (.I(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__A1 (.I(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A2 (.I(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A2 (.I(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__I (.I(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__I (.I(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__A1 (.I(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__A2 (.I(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__A2 (.I(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__I (.I(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A1 (.I(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A1 (.I(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__A1 (.I(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A1 (.I(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__I (.I(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__A1 (.I(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__A2 (.I(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A2 (.I(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A2 (.I(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A2 (.I(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__A1 (.I(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A1 (.I(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__A1 (.I(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__I (.I(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__A1 (.I(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A1 (.I(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__A1 (.I(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06054__I (.I(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__A1 (.I(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__A2 (.I(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A2 (.I(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A3 (.I(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__A2 (.I(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06189__I (.I(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__A1 (.I(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__A2 (.I(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__A2 (.I(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A3 (.I(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__I (.I(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A3 (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A1 (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__A1 (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__A2 (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__A1 (.I(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__A2 (.I(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__A2 (.I(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__A2 (.I(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__A1 (.I(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A1 (.I(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__A1 (.I(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__A1 (.I(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__A2 (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A1 (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__I (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__A1 (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__A1 (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__A1 (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__A2 (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__A2 (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__I (.I(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A2 (.I(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A2 (.I(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A1 (.I(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__A2 (.I(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__I (.I(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A1 (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__A1 (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__I (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__A1 (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__B (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__B2 (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A1 (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__A2 (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__A1 (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__B (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__A1 (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__A2 (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__A1 (.I(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__B (.I(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__A3 (.I(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A1 (.I(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__A1 (.I(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__A1 (.I(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06053__I (.I(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__A2 (.I(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A1 (.I(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__I (.I(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__A1 (.I(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__A1 (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A1 (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A1 (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__A1 (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__B (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__A2 (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__A2 (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__A2 (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A2 (.I(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__A2 (.I(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__A1 (.I(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__A2 (.I(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__A2 (.I(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__B (.I(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__A1 (.I(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__A1 (.I(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__I (.I(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__B2 (.I(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A1 (.I(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A1 (.I(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06061__I (.I(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__A2 (.I(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__A1 (.I(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06243__A1 (.I(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__I (.I(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__A1 (.I(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__A1 (.I(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__C (.I(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__I (.I(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A1 (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__A1 (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__A1 (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__A2 (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__I (.I(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A1 (.I(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__A1 (.I(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__A1 (.I(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__A1 (.I(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__I (.I(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__A2 (.I(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__B (.I(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__B2 (.I(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__A1 (.I(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__A3 (.I(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__A4 (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A1 (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__I (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A1 (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A1 (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__A1 (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__A1 (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06081__I (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06073__B (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__A1 (.I(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06074__I (.I(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A1 (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__B (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__C (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__I (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__I (.I(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__B (.I(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__C (.I(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A2 (.I(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A1 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__A1 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__I (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__A1 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__I (.I(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A1 (.I(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__I (.I(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A3 (.I(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__A1 (.I(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__A1 (.I(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06122__A1 (.I(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__A1 (.I(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__I (.I(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A1 (.I(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__A1 (.I(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A2 (.I(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A1 (.I(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06188__I (.I(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A2 (.I(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__A1 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__A1 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06086__A1 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A2 (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06246__I (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__I (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06086__A2 (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__A2 (.I(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__A2 (.I(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__A2 (.I(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A1 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__A1 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A2 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__A2 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A2 (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A3 (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__I (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__A2 (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A1 (.I(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__A1 (.I(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A1 (.I(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__I (.I(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A1 (.I(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__I (.I(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__A1 (.I(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__A1 (.I(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__A2 (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__A1 (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__A1 (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__A2 (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__C (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__I (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__I (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__I (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__C (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__C (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__I (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__A3 (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__A1 (.I(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__A1 (.I(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A1 (.I(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__A2 (.I(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__I (.I(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__B2 (.I(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A2 (.I(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A2 (.I(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__I (.I(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__A2 (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A1 (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A1 (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06125__A1 (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A1 (.I(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__A2 (.I(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__A1 (.I(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A2 (.I(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A2 (.I(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__A2 (.I(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A1 (.I(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06100__I (.I(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__I (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__A2 (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__A2 (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__A2 (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__I (.I(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06223__I (.I(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__A2 (.I(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A1 (.I(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__A1 (.I(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__A1 (.I(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A1 (.I(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__A1 (.I(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__A2 (.I(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A3 (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__A1 (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A2 (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__A2 (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A1 (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A1 (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__A1 (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__A2 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__A2 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A1 (.I(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A1 (.I(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06125__B (.I(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A2 (.I(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A1 (.I(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A2 (.I(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A2 (.I(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__A3 (.I(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__I (.I(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__I (.I(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A3 (.I(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A2 (.I(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__B2 (.I(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__I (.I(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A1 (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__A3 (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A2 (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A2 (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A3 (.I(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__A4 (.I(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__A1 (.I(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A3 (.I(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A2 (.I(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A3 (.I(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__A3 (.I(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__I (.I(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__B2 (.I(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__A2 (.I(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__A2 (.I(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06160__A1 (.I(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__A1 (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__I (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06136__A1 (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06131__I (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A1 (.I(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A1 (.I(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__A2 (.I(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06134__A1 (.I(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A1 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A2 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__A2 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06134__A2 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__I (.I(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__A2 (.I(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__A2 (.I(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__I (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__I (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__A2 (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__A1 (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A1 (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__I (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A2 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A2 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A3 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__A2 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A2 (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__A2 (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__A2 (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__A1 (.I(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__I (.I(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__A1 (.I(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__A1 (.I(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__A1 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__I (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__I (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__A2 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A4 (.I(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A2 (.I(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__A2 (.I(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A1 (.I(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__A1 (.I(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__A1 (.I(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__I (.I(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A1 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__B2 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__I (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__A1 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A2 (.I(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A2 (.I(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__I (.I(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__A2 (.I(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A1 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__A1 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__B (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__B (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A2 (.I(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__A2 (.I(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__A1 (.I(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__A1 (.I(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__A3 (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__I (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__I (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__A1 (.I(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A3 (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__A3 (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06156__I (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A2 (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A2 (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__A4 (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06157__I (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A1 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__I (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A3 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__A2 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A1 (.I(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__B (.I(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06160__B (.I(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__B (.I(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__A1 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A1 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__A1 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__I (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__A2 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__A1 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__A1 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__B (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A2 (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A1 (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A2 (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__A1 (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__I (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A1 (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A2 (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__I (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A1 (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A3 (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06361__I (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__I (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A2 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A2 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__A2 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06170__I (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__A1 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__A1 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A1 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__I (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A1 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A1 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A2 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__A2 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__A1 (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__A2 (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A3 (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__I (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__I (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A2 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06175__A2 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__I (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A1 (.I(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A1 (.I(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A1 (.I(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__A3 (.I(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A2 (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__B1 (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__B (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__A1 (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__A1 (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06179__I (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__I (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A1 (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__A1 (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__I (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A1 (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A1 (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__B2 (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A1 (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__A1 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A1 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__I (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A2 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__I (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__I (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__B (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A1 (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A3 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__A2 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A4 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__A2 (.I(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__A2 (.I(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A1 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__A1 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A1 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__A1 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__A1 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__A3 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__A2 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__B1 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__C (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__B (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__A1 (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__A1 (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A2 (.I(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A1 (.I(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__B (.I(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A1 (.I(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A1 (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__I (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A2 (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A2 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__I (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A1 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__A1 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__I (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__I (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__I (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A2 (.I(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__A2 (.I(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A2 (.I(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__I (.I(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__C (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__A2 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__I (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A3 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A3 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__A2 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06406__A2 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__A2 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A3 (.I(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__I (.I(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__A4 (.I(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__A1 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A3 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__A2 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__A2 (.I(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11590__A1 (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__A1 (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A1 (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A1 (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__I (.I(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06514__A1 (.I(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__I (.I(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__A2 (.I(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__A2 (.I(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__I (.I(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__I (.I(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__A2 (.I(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__C (.I(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__I (.I(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__I (.I(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A2 (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__I (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__A3 (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A2 (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A3 (.I(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__A2 (.I(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__A1 (.I(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A2 (.I(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__A2 (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__A1 (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__I (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__A3 (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__C (.I(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__A1 (.I(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A2 (.I(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__B1 (.I(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__C (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A1 (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__I (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A2 (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__I (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__B (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__B (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A1 (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__I (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__I (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A2 (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__A2 (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__A2 (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A2 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__I (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__A2 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__A2 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__A2 (.I(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__I (.I(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__I (.I(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__A2 (.I(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A2 (.I(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A2 (.I(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__A3 (.I(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__A3 (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A3 (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__I (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__A2 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A2 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A1 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A1 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__A2 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A2 (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__A2 (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__A2 (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__I (.I(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__B2 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__I (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__I (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__I (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__A2 (.I(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__A1 (.I(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A1 (.I(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__A3 (.I(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__A2 (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__C1 (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__A2 (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__A2 (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__A2 (.I(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__A2 (.I(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__A2 (.I(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__A2 (.I(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A2 (.I(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A1 (.I(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06467__A1 (.I(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A1 (.I(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__I (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A1 (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__A1 (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__I (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__I (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__I (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A2 (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__I (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__A1 (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A1 (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__C (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A2 (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__B (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__I (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__I (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__I (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__A2 (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A2 (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A2 (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06243__A2 (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__A2 (.I(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__A2 (.I(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A1 (.I(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11467__A1 (.I(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__I (.I(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__I (.I(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__A1 (.I(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A1 (.I(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__I (.I(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__A3 (.I(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__A2 (.I(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__A2 (.I(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__I (.I(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A3 (.I(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A2 (.I(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__A2 (.I(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A2 (.I(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A1 (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A1 (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06279__A1 (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__B2 (.I(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A3 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A1 (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__A1 (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__A2 (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__A1 (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__I (.I(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__I (.I(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A1 (.I(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__I (.I(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__C (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11619__C (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11615__C (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A1 (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__A3 (.I(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__A2 (.I(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__A1 (.I(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A2 (.I(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A1 (.I(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06263__I (.I(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A1 (.I(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A1 (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A2 (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A3 (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A1 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__A1 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__A2 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A2 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A1 (.I(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A1 (.I(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__A1 (.I(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A2 (.I(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__A2 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__A1 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__A1 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A2 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__A1 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__I (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__A1 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A3 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__A1 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__A2 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A2 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A3 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__A1 (.I(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__A1 (.I(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__A2 (.I(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__A1 (.I(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__C (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__C (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__I (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__I (.I(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A1 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11476__A1 (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__A2 (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__B (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__I (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__A1 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A2 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__I (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__I (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A1 (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__B (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__I (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__I (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__C (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__C (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__C (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06279__A2 (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__A1 (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A1 (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A2 (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__I (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__A1 (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A1 (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A2 (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__I (.I(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11556__A1 (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A1 (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A2 (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06283__I (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A1 (.I(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A1 (.I(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A1 (.I(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__B2 (.I(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__C (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__C (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A1 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__A1 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__A1 (.I(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__A2 (.I(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__A2 (.I(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A1 (.I(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__I (.I(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__I (.I(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__A1 (.I(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A1 (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__A1 (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__I (.I(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A2 (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__A1 (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06374__A2 (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A2 (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A1 (.I(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__I (.I(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A1 (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A2 (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A2 (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A1 (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__I (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A2 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__A1 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__I (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__I (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__I (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__C (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A3 (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__I (.I(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__I (.I(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__A2 (.I(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__A2 (.I(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A2 (.I(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A2 (.I(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A1 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__B2 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__A1 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__A1 (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__C (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A1 (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__I (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__I (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__I (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__I (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__I (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11617__C (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11585__C (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__I (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__I (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__A1 (.I(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A1 (.I(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__A1 (.I(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A1 (.I(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A2 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A2 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__A2 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__I (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__A2 (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__A1 (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__C (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A4 (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__A2 (.I(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A1 (.I(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A3 (.I(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__A2 (.I(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A1 (.I(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__B (.I(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__A1 (.I(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A2 (.I(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A2 (.I(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A1 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A2 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A2 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A1 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__A1 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__A2 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A3 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A2 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A4 (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A2 (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__A3 (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__I (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A2 (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A2 (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__A2 (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A3 (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__A3 (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A4 (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__B2 (.I(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A1 (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__A2 (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__A1 (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__I (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__I (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__I (.I(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__I (.I(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__I (.I(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__I (.I(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A1 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__A1 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__A1 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__C2 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__I (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__B2 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__I (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__A1 (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A1 (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__A1 (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__I (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__B2 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__I (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A1 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A2 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__I (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__A1 (.I(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__I (.I(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A2 (.I(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A2 (.I(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A1 (.I(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A2 (.I(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__I (.I(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__I (.I(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A2 (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A1 (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A1 (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__I (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__C (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A3 (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__A2 (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__I (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A4 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A2 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A4 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A3 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__A2 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__A2 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__A1 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A2 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A1 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A2 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__I (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__I (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A2 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A1 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A1 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__B3 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__B (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A1 (.I(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A2 (.I(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A2 (.I(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__I (.I(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A1 (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__A1 (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__I (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__I (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__I (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__I (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A1 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__I (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A1 (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A2 (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__A2 (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__A2 (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__B (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__A3 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__I (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__A2 (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__A2 (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A1 (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A1 (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__I (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A2 (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A1 (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__A1 (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__I (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__B2 (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A1 (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A1 (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__I (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A1 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A1 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__A2 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__A1 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A2 (.I(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A2 (.I(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__B1 (.I(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A2 (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__I (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__A1 (.I(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A2 (.I(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A3 (.I(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__A2 (.I(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__C1 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__B1 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__A1 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__I (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__B1 (.I(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__C1 (.I(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__C1 (.I(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__A3 (.I(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A2 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A2 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__A1 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A1 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11507__A1 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__I (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__C (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__I (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A1 (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__A1 (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__B (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A1 (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__B2 (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A1 (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__B (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__A1 (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__A1 (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A1 (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A2 (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A1 (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__A2 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__B2 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__A1 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A2 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A2 (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A2 (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__A2 (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__I (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A2 (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A2 (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A2 (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A2 (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A1 (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__A1 (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__A1 (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A4 (.I(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A1 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A2 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__A2 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A1 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__A1 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A4 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A2 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A2 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__I (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A1 (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A1 (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A2 (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__A2 (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A1 (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A1 (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__A1 (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11570__B2 (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__B (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__A2 (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A2 (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__A2 (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A2 (.I(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__I (.I(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__C (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__I (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__A2 (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__A1 (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A1 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A1 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__A2 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__A1 (.I(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__A2 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__I (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__B (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11227__B (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__I (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__A2 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A1 (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__A2 (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A2 (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__A1 (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__B2 (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__I (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__A3 (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A2 (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__A1 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A1 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__A2 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__A2 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A1 (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A1 (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__I (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A1 (.I(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__B2 (.I(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__A2 (.I(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__A3 (.I(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A3 (.I(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A2 (.I(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A3 (.I(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A2 (.I(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__A1 (.I(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__I (.I(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11544__A2 (.I(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A2 (.I(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A1 (.I(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__A2 (.I(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A1 (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__A1 (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__A1 (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__I (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__A1 (.I(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A1 (.I(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A1 (.I(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__I (.I(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__A1 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A1 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__A1 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__I (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A1 (.I(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__A1 (.I(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__I (.I(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A1 (.I(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A2 (.I(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__A2 (.I(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__B2 (.I(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__A1 (.I(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A3 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A3 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__A2 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A2 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A2 (.I(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__A1 (.I(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06491__A2 (.I(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06427__A2 (.I(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A2 (.I(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__I (.I(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A3 (.I(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__I (.I(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A2 (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A2 (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A2 (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A3 (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A3 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__B (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A1 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__I (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A1 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__I (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A1 (.I(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__A1 (.I(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A1 (.I(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__I (.I(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__A1 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A1 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A1 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__I (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__C (.I(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__C (.I(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__C (.I(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A1 (.I(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A3 (.I(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A1 (.I(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A4 (.I(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A2 (.I(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__A1 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A1 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__A1 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__I (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A1 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__A1 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A1 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__I (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A1 (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A2 (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A1 (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A1 (.I(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A2 (.I(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A4 (.I(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__B1 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__A1 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__B2 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06446__A1 (.I(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__B (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A2 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A2 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__I (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A1 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__I (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__A3 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06449__I (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A2 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__A2 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__A1 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06450__I (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__A2 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__A2 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__A1 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A2 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A1 (.I(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__A2 (.I(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A2 (.I(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A2 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A1 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__A2 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__B2 (.I(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__A2 (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A1 (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A1 (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__B1 (.I(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A2 (.I(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A2 (.I(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__A1 (.I(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A2 (.I(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A2 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A1 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A4 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__A4 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__B2 (.I(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__C (.I(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A1 (.I(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A2 (.I(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__A1 (.I(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__B (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__B (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__B (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__B (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__B1 (.I(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__A2 (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__C (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A2 (.I(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A1 (.I(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A1 (.I(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__A1 (.I(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__A2 (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__I (.I(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A2 (.I(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__I (.I(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A2 (.I(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A3 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A2 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A2 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__A2 (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A3 (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A3 (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__A1 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__I (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A1 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__A1 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__A1 (.I(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__I (.I(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A2 (.I(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__A2 (.I(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__A1 (.I(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A1 (.I(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__A2 (.I(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__A2 (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__I (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06489__I (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__A2 (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__A2 (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A2 (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__A1 (.I(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__A2 (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06493__I (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A2 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__I (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__A2 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A2 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A1 (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__B2 (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__A1 (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__A2 (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A1 (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A1 (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A2 (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__A2 (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__C (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__C (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__I (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__I (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__C (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__B (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__A2 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A2 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__I (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__I (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06503__A2 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A1 (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__A1 (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__A2 (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__A1 (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__I (.I(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__A1 (.I(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A1 (.I(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__A1 (.I(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11556__A3 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__A2 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__I (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__A2 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__A2 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__B2 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__A1 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__B1 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A1 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A2 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__A2 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__A1 (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A1 (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__I (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A1 (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A4 (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__B (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__I (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__I (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__I (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__I (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A3 (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A2 (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A1 (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__A1 (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__A2 (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A1 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__I (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A2 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A2 (.I(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A2 (.I(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__A2 (.I(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__A3 (.I(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A1 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A3 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__A1 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__I (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A2 (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A1 (.I(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__B (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A2 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A2 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__A2 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__S (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__I (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__I (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A3 (.I(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A1 (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__C (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A2 (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A2 (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A2 (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__I (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A3 (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A1 (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__A2 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A2 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__A4 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A2 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__A2 (.I(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A2 (.I(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A2 (.I(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__A2 (.I(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A2 (.I(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__I (.I(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A1 (.I(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A1 (.I(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__A1 (.I(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A2 (.I(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__A2 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__A2 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__A2 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__A2 (.I(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__I (.I(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A3 (.I(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08825__A1 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A2 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06540__A2 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__I (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A2 (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A3 (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__A3 (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08825__A2 (.I(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A3 (.I(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06540__A3 (.I(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A3 (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A2 (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__A3 (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__A3 (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__A1 (.I(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A2 (.I(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__A2 (.I(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__A2 (.I(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A2 (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__I (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__I (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__I (.I(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A2 (.I(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__A2 (.I(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__A2 (.I(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__I (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A1 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A1 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A1 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__A2 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A3 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__A3 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__A3 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A1 (.I(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__C (.I(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__A1 (.I(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__A4 (.I(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__A2 (.I(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__A2 (.I(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A1 (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A1 (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__A1 (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A1 (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A1 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06607__A1 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A1 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A1 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__I (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__B (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__B (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A4 (.I(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A3 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__A2 (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__A2 (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A4 (.I(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__C (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__A1 (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A2 (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A2 (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__I (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A2 (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06567__I (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A2 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__A2 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A2 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__A2 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__A1 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__B (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__A1 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__I (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A1 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__A1 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A1 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A2 (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A2 (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__A2 (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__A2 (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A3 (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__I (.I(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A1 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__A2 (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__A1 (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__B2 (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__A1 (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__I (.I(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__A3 (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A2 (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__B (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__I (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__A1 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A1 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__I (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__A1 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A2 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A3 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__A2 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__A2 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__A2 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A1 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__A1 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A1 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A2 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__C (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__B (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__I (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__A1 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__A1 (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__I (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A1 (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A1 (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A1 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A1 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__A1 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A2 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__I (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__B2 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__I (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__A2 (.I(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__B (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__B (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__B (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__A2 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A1 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A2 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__A2 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__A1 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__I (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A2 (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__I (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__A1 (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__B (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__B (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__I (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__I (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__I (.I(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A3 (.I(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A2 (.I(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A2 (.I(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__B (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__B2 (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__A2 (.I(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A1 (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__A1 (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A2 (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06598__I (.I(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__B2 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__B1 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__A2 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__I (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__A1 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A1 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06607__A2 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__C (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__I (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__I (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__B (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__C (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A2 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__B (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__A3 (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__A1 (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__C (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__C (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__B (.I(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A2 (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__A1 (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__B (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__B2 (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__I (.I(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__A1 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__A1 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__A1 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__A1 (.I(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A1 (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__A1 (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__I1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__A1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__A1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__A1 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__I (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__C (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__A2 (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__C (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__A2 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A3 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__A1 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__A3 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__I (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__B1 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__B (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__A1 (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__I (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__B2 (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A1 (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A2 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__A1 (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__I (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__A1 (.I(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A1 (.I(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__B2 (.I(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__A1 (.I(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__I (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__A1 (.I(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__A2 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06644__I (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07059__I (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__B2 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__B2 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__B2 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__A2 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A2 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__A1 (.I(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__A1 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A1 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A2 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__A2 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__B2 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__A1 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A3 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__A3 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__B2 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__A1 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A1 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__C (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A1 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A1 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__A1 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__B2 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A2 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A1 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__A2 (.I(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__I (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A2 (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A1 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__A1 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07368__A1 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06657__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__A1 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__B2 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__I (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__I1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A1 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A1 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__I (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A1 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A2 (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A3 (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A3 (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A3 (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__A1 (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__I (.I(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__A2 (.I(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__I (.I(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__A2 (.I(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__I (.I(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__A2 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__I (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__A2 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__A2 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__A2 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__I (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A2 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__A2 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A3 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__I (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A2 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__A1 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__A2 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__A3 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A2 (.I(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__A2 (.I(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__A2 (.I(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__A2 (.I(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09642__A2 (.I(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A2 (.I(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__I (.I(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__A1 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__A1 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__I (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__A1 (.I(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__A2 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__A2 (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__B (.I(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__A2 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__I1 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__A2 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__I (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A3 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__A3 (.I(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__C (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__I (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A4 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A3 (.I(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A2 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__A3 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A2 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__A3 (.I(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__B (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__I (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__I (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__A2 (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A1 (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__B (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__I (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A1 (.I(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A1 (.I(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__I (.I(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A1 (.I(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11433__A1 (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__A2 (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07032__A2 (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A2 (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__B1 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A1 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A1 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__I (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__B2 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__A2 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A1 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A2 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__I (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__A1 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__B1 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__I (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A1 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A1 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A1 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__A1 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__B (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__B (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__I (.I(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__A1 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__A1 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__A1 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__B1 (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__A1 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__A1 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__A1 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A1 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__A2 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A2 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A1 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__I (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__A2 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A2 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A2 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__B (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A3 (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__A2 (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A2 (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__A2 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A1 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__A2 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__C (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__C (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__C (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__I (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__A1 (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07060__C (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A1 (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__A1 (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__A1 (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A1 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__A2 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__A3 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__B1 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A1 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__A1 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__A1 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__A1 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A2 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__A2 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__A2 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A1 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__A2 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A1 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A2 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__I1 (.I(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__I (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__A2 (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A2 (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__A2 (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__I (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__I (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__A1 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07413__A1 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__A1 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A2 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A2 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__A1 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__B1 (.I(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__A1 (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__B1 (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__A1 (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__I (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__B (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__A1 (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A2 (.I(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__A4 (.I(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__B1 (.I(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__A4 (.I(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A2 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__I (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__I (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A1 (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__A2 (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__A2 (.I(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__A2 (.I(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__A2 (.I(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A1 (.I(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__B1 (.I(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A1 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__A1 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__B2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__B2 (.I(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__B (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__B (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__I (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__A1 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__B1 (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__A1 (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__A1 (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A2 (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__B (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__B (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__I (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__I (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A2 (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__A1 (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__A1 (.I(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__B2 (.I(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__A2 (.I(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__A2 (.I(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__C (.I(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A2 (.I(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__B1 (.I(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__A2 (.I(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__A2 (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A2 (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__A2 (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A2 (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A3 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__A2 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__C (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__I (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__I (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__A2 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A1 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__A1 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A3 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__A3 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__A2 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A1 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A1 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__A1 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A1 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__A2 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A2 (.I(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__A1 (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__A1 (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__B (.I(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__A3 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A2 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A2 (.I(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__A4 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A3 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A3 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__A2 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A2 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__I1 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__A2 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11533__A1 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A1 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A1 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__I (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__I (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A1 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A1 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__A1 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A4 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A1 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__I (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A1 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__A1 (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A2 (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A1 (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__I (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A1 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__A1 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__A1 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__A1 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A1 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__A2 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08575__I (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__I (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__A1 (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A1 (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A1 (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A1 (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__A1 (.I(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A1 (.I(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A1 (.I(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A2 (.I(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A2 (.I(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__A2 (.I(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__A2 (.I(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A4 (.I(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A3 (.I(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A3 (.I(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A2 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A2 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A1 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__A2 (.I(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11609__A1 (.I(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A1 (.I(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A1 (.I(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A1 (.I(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__I (.I(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__C (.I(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__C (.I(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A2 (.I(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11433__A4 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__I (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__A1 (.I(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A1 (.I(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__A2 (.I(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__A2 (.I(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A1 (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__B1 (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__I (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__A1 (.I(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A2 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A2 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__B1 (.I(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__B2 (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__B2 (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__A1 (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__B2 (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A2 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__A2 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__I (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A2 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A2 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A1 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__A2 (.I(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A4 (.I(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__B (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A1 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__A1 (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A1 (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__I (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A1 (.I(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__I (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A1 (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__A1 (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A1 (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A2 (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__I (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A2 (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__A1 (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A2 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__A1 (.I(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__A1 (.I(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A1 (.I(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A1 (.I(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__B2 (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__B2 (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__I (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__B2 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07156__A1 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__B2 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A1 (.I(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A2 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__B1 (.I(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__A2 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__A2 (.I(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11567__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07150__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06908__A1 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__I (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A1 (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__B2 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__A2 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__A2 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A2 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07149__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07060__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__A1 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__B1 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__A1 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__A1 (.I(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A2 (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A2 (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__B (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__B (.I(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__A2 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A1 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A4 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__I1 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__I (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A2 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__B2 (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__A1 (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06936__A1 (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__A1 (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A2 (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A2 (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__I (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A3 (.I(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__B (.I(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A2 (.I(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__A1 (.I(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__I (.I(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A2 (.I(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A1 (.I(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__B1 (.I(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__A1 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__B1 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__A2 (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06939__I (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A2 (.I(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__I (.I(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__B1 (.I(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__A2 (.I(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07067__A2 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A2 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__B1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__I (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__A1 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__A1 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__A1 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06974__A1 (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__A1 (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__A1 (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__A1 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__A1 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__I (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__A1 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__I (.I(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__A2 (.I(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A2 (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__B (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__A2 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__C (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__B2 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A3 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__A3 (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__A1 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__A1 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__B1 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__A3 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__I (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__A2 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__I1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A2 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A2 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__A2 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__B1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__B1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__A2 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A2 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__I (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__A2 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A2 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A1 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__A2 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A3 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07495__I (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__A1 (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A1 (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A1 (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__I (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A2 (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__I (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__A1 (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__A1 (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A2 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__C2 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__B1 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__I (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__I (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__B1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__I (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A1 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__A2 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__A2 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__A2 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A1 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07010__A2 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__A2 (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__A1 (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__I (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A1 (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A1 (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__A2 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__B1 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A3 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A2 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__A2 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A1 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__B1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__C1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__I (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A2 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A2 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__I1 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A2 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A2 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__I (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07032__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__C1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__A3 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__I (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11584__A1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__A1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__B1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__A2 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__I (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__I (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__I (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A1 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A1 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__B1 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A1 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__C (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A2 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A2 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__A2 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__I (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__A2 (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A2 (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A1 (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__A2 (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__I1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__B1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07144__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A2 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__B (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A3 (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07058__A1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__A1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A2 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A2 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A2 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__A2 (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A2 (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__B2 (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07060__B2 (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__A2 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__A2 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__I1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__I (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A2 (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A2 (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__A2 (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07077__I (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A2 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A2 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A3 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07079__I (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A2 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A2 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A1 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__A2 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__A1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07088__A1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__A2 (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07088__A2 (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__B1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__A2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__I (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__A1 (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A1 (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07114__A1 (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__A1 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__A1 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__A2 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__B1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__I (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__A1 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A1 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A1 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__I (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__B (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11566__A2 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A2 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__A2 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11291__A2 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__A3 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__A2 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__B1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__A2 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__C1 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07156__A2 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A2 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A1 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__A2 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__I (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A1 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A1 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__I (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A1 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__A1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__A1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A2 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__I (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__I (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A1 (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A2 (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A2 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A2 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__I (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__A1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A2 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A2 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07177__A2 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A2 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__I (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__A2 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__A2 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__A2 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__A1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__A2 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__A1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__A1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A3 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__A1 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A2 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__I (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__A3 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__A2 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A1 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__B1 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A1 (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A1 (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__I (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__I (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__I (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__A1 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A1 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A2 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A1 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__S (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A2 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__I (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A1 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A2 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__A2 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__A2 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__B2 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A2 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__B1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__B1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__A2 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__A2 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__A2 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A2 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__I (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A2 (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A2 (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__I (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__A2 (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__A2 (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__A1 (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__A2 (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A1 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__I (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__I (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__A1 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__B1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A2 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A2 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__A2 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__A1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__A1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__A2 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__I (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__A2 (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__A2 (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A2 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A3 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A2 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A4 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A2 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__I (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__I (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__A3 (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A2 (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__I (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A2 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07732__A2 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__I (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__A2 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A2 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__A1 (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__B (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A1 (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__I (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__A1 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__I (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__I (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__I (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__B (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__B (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A1 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__A1 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__A2 (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__I (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__A1 (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__I (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__A2 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__A2 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07404__I (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__I (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__I (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__I (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__A2 (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__I (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__C2 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__A2 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__A2 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__A2 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10569__I (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__B1 (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__B1 (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__I (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__B1 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__B1 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A2 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__I (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__I (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__I (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A2 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__I (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__I (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__C2 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A2 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__B1 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__B1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__A2 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__B1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07316__I (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__B1 (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__B1 (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__B1 (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07320__I (.I(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__B1 (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__B1 (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__B1 (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__I (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__B1 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__B1 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__I (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__I (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__B1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__B1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__B1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__B1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__I (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__B1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__B1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__B1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__I (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__B1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__A2 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__C1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A1 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A1 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__B (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__I (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__A1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__A1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07348__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07330__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__B (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__A2 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__I (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__A2 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A1 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A1 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A1 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__A1 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__B2 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__I (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__A1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A2 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__A2 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11542__A1 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07557__I (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__A2 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__B (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__A1 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__I (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07340__I (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__B (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__A1 (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A1 (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__I (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__I (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__B (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__I (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__B (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__B1 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__A2 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__B1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__B1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__I (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__A2 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__A2 (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__I (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__I (.I(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__I (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__I (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A2 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__C2 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__A1 (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A1 (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A1 (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__B (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__B (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__B (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__A1 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__I (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__A1 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A1 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A1 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07352__I (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__I (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__B (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__B (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__A1 (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__B1 (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A2 (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A2 (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__I (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A2 (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__B1 (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__A2 (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__I (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__I (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__I (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__I (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__B1 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__B1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__B1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__B1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__I (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__B1 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__B1 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__B1 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__I (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__I (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__I (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__I (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__B1 (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__B1 (.I(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__A2 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A1 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__A2 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__A1 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__A1 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A2 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A2 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__I (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__I (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__A2 (.I(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__I (.I(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__I (.I(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__I (.I(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__I (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__I (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__I (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__I (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__A2 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__A2 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__B1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__A2 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__A2 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__B1 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__I (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__I (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__I (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__I (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__B1 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A2 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__A2 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__B1 (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__B1 (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__B1 (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__I (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__B1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__B1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07445__I (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__I (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__I (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__I (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__B1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__B1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__B1 (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__B1 (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__I (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07388__I (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__B1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__B1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A2 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__I (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__I (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__I (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__I (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__A2 (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__B1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__B1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__B1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__I (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__B1 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__B1 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__B1 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07392__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__B1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__B1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__A2 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__A2 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__B1 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__I (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__A2 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__A2 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__A2 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__I (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__I (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__I (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__A2 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__C1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__I (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A2 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A2 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__A2 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A2 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__A2 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__A2 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__I (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A2 (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__A2 (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__A2 (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A2 (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__B (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__A1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__B2 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__B (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__I (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__B2 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A1 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__B2 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__I (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__B (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__B (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__B (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__B2 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__I (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A2 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A1 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A1 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__A1 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A1 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__I (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__B1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A2 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A2 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__B1 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__B1 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__B1 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__B1 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A2 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A2 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__A2 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__A2 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__A2 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__C1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__B1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__B1 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__A1 (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A2 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A2 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A2 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11207__I (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__B1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__B1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__B1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A1 (.I(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A2 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A2 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A2 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__A2 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__B (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__B (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__B (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__B (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__I (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__A2 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A2 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A2 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__I (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__I (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__C2 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__C2 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__B (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__B (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__B (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__B (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__I (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__A2 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__A2 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A2 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__C2 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__C2 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A2 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__I (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11508__A2 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__C2 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__C2 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__I (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__I (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A2 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__B1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__B1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11214__I (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__B1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__B1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__B1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A3 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__B (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__B1 (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__A1 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A1 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07452__A2 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__A1 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A1 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A1 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__I (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__I (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__B1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A2 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A3 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__B (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__B1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A1 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A1 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A2 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__I (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__A1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__A1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__A2 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__A2 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A2 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__A2 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__C2 (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__I (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A2 (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__A2 (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__B1 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A2 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__I (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A2 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A1 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__B (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__B1 (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A1 (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A1 (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A2 (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__A1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__I (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A1 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__B (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__C2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A1 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A2 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__A2 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__A1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__B1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__B1 (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__B1 (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__B1 (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__A2 (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__C1 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__B1 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__I (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__B1 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__A2 (.I(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__I (.I(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__C2 (.I(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A2 (.I(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__I (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__B1 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__B1 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__B1 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__B1 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__I (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A2 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__C1 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__A2 (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__B1 (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__A2 (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__A2 (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A2 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__B (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A1 (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A1 (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A2 (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__I (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__C2 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__A2 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A2 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__A2 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__B1 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__B1 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__B1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__B1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__B1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__B1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__B (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__B1 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__A1 (.I(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__A1 (.I(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__A2 (.I(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__I (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__A1 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A1 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A1 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__B (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A1 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A1 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A1 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__A1 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__B (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__A1 (.I(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__I (.I(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__I (.I(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__I (.I(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A1 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A1 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07740__A1 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A1 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A1 (.I(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A1 (.I(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A1 (.I(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07568__A1 (.I(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__A1 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11510__A1 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__B1 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__A3 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__I (.I(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__I (.I(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__I (.I(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__I (.I(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07568__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A1 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A1 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__I (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__A1 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__A1 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__A1 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A1 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__I (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__I (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07716__A2 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__I (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__A2 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07618__I (.I(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__I (.I(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__A2 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__A2 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A2 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A2 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A1 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A2 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A2 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__I (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__I1 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A2 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A2 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A2 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__A2 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__B1 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__B1 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__I (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__A1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__A1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A3 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A2 (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__A2 (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A2 (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__A1 (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A2 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__A2 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__A2 (.I(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__A2 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__I (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__I (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__B2 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__A3 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__I (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A1 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__I (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__A2 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__A2 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__I (.I(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__B (.I(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__A2 (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__A2 (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__I (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__A2 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A2 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A4 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A4 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A4 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A4 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__I (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__I (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__A2 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__A2 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__A2 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__A2 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11550__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11547__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__A1 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__B2 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__A1 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A2 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__I (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__I (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__A1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__I (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08155__I (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__I (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__I (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A3 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A3 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__A3 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A3 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__I (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__I (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__I (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__I (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__A1 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A1 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__I (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__I (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__A3 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__I0 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__I0 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__I (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__A2 (.I(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__A2 (.I(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__I (.I(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A1 (.I(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__I (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__I (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__I (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__I (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__A1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__A2 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__I (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__I (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__I (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__I (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__C (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__C (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__C (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__B (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__I (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A1 (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__I (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11619__A1 (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__I (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__I (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__I (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A1 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A1 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__A1 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A1 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__A2 (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__A1 (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__I (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__I (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__A1 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__A1 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__A1 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__A1 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A2 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__B1 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__A2 (.I(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A2 (.I(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__A2 (.I(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A2 (.I(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__B (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__B (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__B (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__B (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A1 (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__I (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__I (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__I (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__I (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__I (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__A1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__A1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__A1 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__B (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__A1 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__I (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__A1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__A1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__I (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__I (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__I (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__I (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__A1 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A1 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A1 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__A2 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__B2 (.I(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__A1 (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__I (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__C1 (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__I (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11615__A1 (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__I (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__I (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__I (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A1 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A1 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A1 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__A1 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__A3 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__I (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A1 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__I (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__A1 (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A1 (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__I (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A1 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__B (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A1 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A1 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__I (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__I (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__I (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__I (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A1 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A1 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A1 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A2 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__B2 (.I(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A1 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A1 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__B2 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__I (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__I (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__I (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__I (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__I (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A1 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A1 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A1 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A1 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A2 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A2 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A2 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A2 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__A1 (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A1 (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__I (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A1 (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__A1 (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__A1 (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__I (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__I (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__I (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__I (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A1 (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A1 (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__A1 (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__A2 (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__I (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__B2 (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__I (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11587__A1 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__I (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__I (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__I (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__A1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A2 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A1 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A1 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__A1 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__A1 (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__B2 (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__A1 (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__I (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__A1 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__B (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__A1 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__A1 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__I (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__I (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__I (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__I (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__A1 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A1 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A1 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__A2 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__B2 (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__I (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__I (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__I (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__I (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A1 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__A1 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A1 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A1 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__A1 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A1 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__I (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__I (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A1 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__A1 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__A1 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__I (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__I (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__I (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__I (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__A1 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A1 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A1 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A2 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__B2 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__I (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__I (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__I (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__I (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A1 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A1 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__A1 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__I (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A1 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__B2 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A1 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A1 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__I (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__I (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__I (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__I (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__A1 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__A1 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A1 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A2 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__I (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__I (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A1 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A1 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A1 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A1 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__A1 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A1 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__I (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07716__A1 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A2 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A2 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__I (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__A2 (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A2 (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A1 (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A3 (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__I (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__I (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__B (.I(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__B (.I(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__B (.I(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__I (.I(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A2 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__A2 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__A2 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__I (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A1 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A1 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A3 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A1 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__A2 (.I(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__A2 (.I(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A2 (.I(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A3 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A3 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__A3 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A3 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__I (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__I (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A2 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A2 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__A2 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A2 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__A1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11542__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A1 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__I (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__A1 (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A1 (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A1 (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__A1 (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__I (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__I (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__I (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__I (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__I (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__I (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__I (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__I (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__C (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__C (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__C (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__B (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__A2 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A2 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__I (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__I (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A1 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__A1 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A1 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A2 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A2 (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07766__A2 (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A2 (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__A2 (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__A1 (.I(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A1 (.I(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A1 (.I(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__A1 (.I(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A1 (.I(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A1 (.I(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A1 (.I(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A1 (.I(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__A2 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A2 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A2 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A2 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07908__A1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__A1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A1 (.I(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A1 (.I(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A1 (.I(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A1 (.I(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A2 (.I(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A2 (.I(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__A2 (.I(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A2 (.I(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__A1 (.I(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A1 (.I(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A1 (.I(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__A1 (.I(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__A1 (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A1 (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__A1 (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A1 (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A1 (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__A1 (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A1 (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A1 (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__I (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__I (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__I (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__I (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A1 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A1 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A1 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A1 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A1 (.I(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__A1 (.I(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__A1 (.I(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__B2 (.I(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__I (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__I (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__I (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__I (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A2 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__A1 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A2 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A2 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__I (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__I (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__I (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__I (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__I (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__I (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__B (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__C (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__C (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__B (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A2 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A2 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A2 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A2 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__A1 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__A1 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__A1 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__B2 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A2 (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A1 (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__A2 (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A2 (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A2 (.I(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__A2 (.I(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__A2 (.I(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__A2 (.I(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__C (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__C (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__C (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__C (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A1 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A1 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A1 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__B2 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__I (.I(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__I (.I(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__I (.I(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__I (.I(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A2 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__A1 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A2 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A2 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__A1 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A2 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A1 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__I (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A1 (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A1 (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A1 (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__B2 (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__I (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__I (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__I (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__I (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A2 (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__A1 (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__A2 (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A2 (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A2 (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__A1 (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A1 (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__A1 (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A2 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A2 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__B1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__A1 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__A1 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__A1 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__B2 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A2 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__A2 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__A2 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__B2 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__I (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__I (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__I (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__I (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__A2 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A2 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A2 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__A2 (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A2 (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A2 (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__I (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__B2 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__A2 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A2 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A1 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__I (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__B2 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__I (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__I (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__I (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__I (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A2 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A1 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A2 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__A2 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__A1 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A1 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__A1 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A1 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__A2 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A2 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A2 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A2 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A1 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A3 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__I (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__I (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__I (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__I (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__A2 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__A2 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A2 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__A2 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A3 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A3 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A3 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A3 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__I (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__I (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__I (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__I (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__I (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__I (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__B (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__B (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__B (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__C (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A2 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__A2 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A2 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__A2 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A2 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__A2 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__A2 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A2 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__A2 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A2 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A2 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__A2 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__B (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__B (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__B (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__B (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__B (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__B (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__B (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__I (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11346__A2 (.I(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__B1 (.I(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__B1 (.I(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__I (.I(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A3 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A2 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__A2 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A2 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A2 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__A1 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A1 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A1 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A1 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__I (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__I (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__I (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__I (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__A2 (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__A2 (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__I (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__I (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A2 (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07958__A2 (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A2 (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A2 (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__I (.I(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__I (.I(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__I (.I(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__I (.I(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__C (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07958__C (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__C (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__B (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__B2 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A1 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__A1 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A1 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__A1 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A2 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__A2 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__A2 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A2 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A2 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A2 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A2 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A2 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__B2 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A2 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A2 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A2 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A2 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__C (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__C (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__C (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__C (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__B (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__A1 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A1 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A1 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__A1 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A2 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A2 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A2 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A2 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__A1 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A1 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A1 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A1 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__A1 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__A1 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A1 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A1 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__A1 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A1 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A1 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07958__A1 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__B (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__B (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__I (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__I (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A2 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A2 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A4 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__I (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__C (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__C (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__C (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A1 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__A3 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A2 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A2 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A3 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A2 (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__I (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A4 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__B (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__A1 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A2 (.I(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A2 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__I (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__A1 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A1 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A1 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A1 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A1 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A1 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__I (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09271__A1 (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A1 (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A1 (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__I (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A2 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__I (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__I (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__B (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A1 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__I (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__I (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11533__C (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__C (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__I (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__I (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__B (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__I (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A1 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A2 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__C (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A2 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__B (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__B1 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__B (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__B (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__B (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__I (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A2 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A2 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A2 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A2 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__I (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__I (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A2 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A2 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A2 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A2 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A2 (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A2 (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A2 (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__A2 (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__A1 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A1 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A1 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A1 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__B (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__B (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__B (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__B (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A2 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A2 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A2 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A2 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__A1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__C2 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__A2 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__C2 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__I (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A3 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A2 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A2 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A2 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A2 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__B2 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A1 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__A1 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A1 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__A1 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__B1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A1 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A1 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A1 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__A1 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__A1 (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__A1 (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__A1 (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A1 (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A2 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__A2 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A2 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A2 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A1 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A1 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A1 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A1 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A1 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__A1 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A1 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__A1 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A1 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__A1 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A1 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A1 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__I (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__I (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__I (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__I (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A2 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__I (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A2 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__I (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A2 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A2 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A2 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A2 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__I (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__I (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__I (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__I (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__B (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__B (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__B (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__C (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A2 (.I(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A2 (.I(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A2 (.I(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A2 (.I(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A2 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A2 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A2 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A2 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A2 (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A2 (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A2 (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A2 (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__B (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__B (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__B (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__B (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__B (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__B (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__B (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__I (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A2 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A2 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A2 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__A2 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__A2 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A2 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A2 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A2 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__B (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__B (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__B (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__B (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A1 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A1 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A1 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A1 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A2 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A2 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A2 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__A2 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__I (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__I (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__I (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__I (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A2 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A2 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A2 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A2 (.I(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__I (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__I (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A3 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A3 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A3 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A3 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__I (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__I (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__I (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__I (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__B (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__B (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__B (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__C (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__A2 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A2 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A2 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__A2 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__B (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__B (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__B (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__B (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A2 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__I (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A2 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__I (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__A2 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A2 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__A2 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A2 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A2 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A2 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A2 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A2 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__I (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__I (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__I (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__I (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__I (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__I (.I(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__B (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__B (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__B (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__C (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A2 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A2 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A2 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A2 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A2 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__A2 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A2 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__A2 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__B (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__B (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__B (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__B (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__I (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__I (.I(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__A1 (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__A2 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A2 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A2 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__A2 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A1 (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__A1 (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__A1 (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A1 (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__A1 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A1 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A1 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A1 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A1 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A1 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__A1 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A1 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A1 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A1 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A1 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__A1 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08212__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__I (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__I (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__I (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__I (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__I (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__I (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__I (.I(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__I (.I(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__I (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__I (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__I (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__I (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A2 (.I(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A2 (.I(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A2 (.I(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A2 (.I(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A2 (.I(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A2 (.I(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__A2 (.I(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A2 (.I(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A2 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A2 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A2 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__I (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__A3 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A2 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A3 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__B (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A2 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A4 (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A3 (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__A3 (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A4 (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A1 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A1 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A1 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A1 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A2 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__I (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A4 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A2 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A4 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A4 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A2 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A1 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A3 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__I (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__I (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__I (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A4 (.I(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A1 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__B (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A1 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A1 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A2 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__A1 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A2 (.I(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__B1 (.I(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__I (.I(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A1 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A2 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A1 (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__I (.I(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11603__A2 (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A1 (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__A2 (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__A2 (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__B (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__A2 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A2 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__I (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__I (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A3 (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A2 (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__A2 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A3 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__A2 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A4 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A4 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__A1 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A2 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A2 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__C (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A3 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A4 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A2 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__I (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A1 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A1 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A1 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A2 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__I (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A2 (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__A2 (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__A1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A2 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__C (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__A2 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A1 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__B (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__B (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__A2 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__A1 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__I (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__I (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A1 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A2 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A2 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__B2 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A2 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A2 (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A3 (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A1 (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A1 (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__I (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__A1 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A3 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A3 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A3 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__A3 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__A2 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A2 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A1 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A2 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A1 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A3 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__A1 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A3 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A2 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__A2 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__B2 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__C (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__I (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__I (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11581__A2 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__B (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__A1 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A1 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__B2 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A1 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A1 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__A2 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__A1 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A1 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__I (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__A1 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A1 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A2 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__I (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A1 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11627__A1 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11623__A1 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__I (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A2 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11521__A1 (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A1 (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A2 (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__I (.I(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10607__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__C (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__B2 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__B2 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__A1 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__B (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__C (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__I (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__I (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__I (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__I (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__I (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__I (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A2 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A2 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__I (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__I (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__I (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__I (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__I (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__I (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__B (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__B (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__B (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__C (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A2 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__A2 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A2 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__A2 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__A2 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__A2 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A2 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__A2 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__B (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__B (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__B (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__B (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__I (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__I (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__I (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__I (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A2 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__I (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A2 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__I (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11540__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A2 (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A2 (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A2 (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A2 (.I(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09344__I (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08350__I (.I(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__B (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__B (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__B (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__C (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__A2 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A2 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A2 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A2 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A2 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A2 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A2 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A2 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__A1 (.I(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A1 (.I(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A1 (.I(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A1 (.I(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__A3 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__A3 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A3 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A3 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09289__I (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__I (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__I (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__I (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A2 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A2 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A2 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A2 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__I (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__I (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__I (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__I (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__B (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__B (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__B (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__C (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__A1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__A1 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__A1 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A1 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A1 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__A1 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A1 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A1 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__A1 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__A2 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A2 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A2 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__A2 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__B (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__B (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__B (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__B (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A1 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08448__A1 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A1 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A1 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__I (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__I (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__I (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__I (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__A2 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__I (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A2 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__I (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A2 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A2 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A2 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A2 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__I (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__I (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__I (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__I (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__B (.I(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__B (.I(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__B (.I(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__C (.I(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A2 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A2 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__A2 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A2 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__B (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__B (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__B (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__B (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__I (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__I (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__I (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__I (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__I (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__I (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__B (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__B (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__B (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__C (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__A2 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__A2 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A2 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A2 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A2 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08448__A2 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A2 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A2 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__B (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08448__B (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__B (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__B (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A2 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__I (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A2 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__I (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__A2 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__B (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A1 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__A1 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A1 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__A1 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__B (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__A3 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__A2 (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__A1 (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A2 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A2 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A3 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A3 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11554__A2 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A2 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__A2 (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A1 (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A1 (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11563__A3 (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A1 (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A2 (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11556__A4 (.I(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A3 (.I(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11603__A1 (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A2 (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A3 (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__A1 (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A3 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__B1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__B2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__C (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__A3 (.I(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A2 (.I(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A2 (.I(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A4 (.I(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__B (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A2 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A1 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__I (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A1 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A1 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__I (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__A2 (.I(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A2 (.I(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A1 (.I(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A2 (.I(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A1 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__B (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__B (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A2 (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11563__A2 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A2 (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__A2 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__I (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__B1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A2 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A3 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A2 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__A1 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A4 (.I(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A2 (.I(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__B (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A2 (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A1 (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__I (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__I (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A1 (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__A3 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A4 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__A2 (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__I (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__I (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A3 (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__A4 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A3 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A2 (.I(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__B (.I(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__A1 (.I(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A2 (.I(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11531__I (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__A1 (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__I (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__I (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__A1 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__A1 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A1 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A1 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__B2 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__A1 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__A1 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A1 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__I (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__I (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__B1 (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A2 (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A2 (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A2 (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__A1 (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10575__A1 (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A1 (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A1 (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A1 (.I(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__B1 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__B1 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__I (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__I (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__B1 (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__B1 (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__B1 (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__B1 (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__A2 (.I(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__C2 (.I(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__C2 (.I(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__A2 (.I(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A2 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A2 (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__A2 (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A2 (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__A1 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__B (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A1 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__A1 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__B (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__A1 (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A1 (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__I (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__I (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__A2 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A1 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__I (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A2 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A1 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A2 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__I (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__C (.I(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A1 (.I(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A1 (.I(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A1 (.I(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__A1 (.I(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__A3 (.I(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A1 (.I(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__A1 (.I(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__A2 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A1 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__A2 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A1 (.I(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A2 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__B (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__A1 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__I (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__A2 (.I(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__A2 (.I(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__A2 (.I(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__A2 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__C (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__A1 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__A1 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A3 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__B (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A1 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__I (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__I (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__I (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__C (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__I (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__I (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__C (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__I (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__I (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A2 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A2 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__A3 (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11584__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A1 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__A1 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__A1 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__A1 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__A1 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__B2 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A1 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__A2 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A1 (.I(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__A1 (.I(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__B1 (.I(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__I (.I(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__A1 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A1 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__A1 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__A4 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A3 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11556__A2 (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A1 (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__A1 (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__I (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A1 (.I(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A3 (.I(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A1 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__I (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__A1 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A2 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__I0 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A1 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__A1 (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__A1 (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A1 (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__I (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__A1 (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__I (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A2 (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A2 (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A1 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A1 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A2 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__I (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A2 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__I (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__I (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A2 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A1 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__I (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__B2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__A1 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__A1 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A3 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A1 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A1 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A1 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__I (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A1 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__A1 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__B2 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__I (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__C2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__I (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__A1 (.I(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__I (.I(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__A1 (.I(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__I (.I(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__A1 (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__B2 (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__A1 (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A4 (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__A1 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__A2 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A1 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__I (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__I (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A3 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__A1 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__B2 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A1 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__A1 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__I (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__A1 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A3 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__I (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A2 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A2 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A2 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__A2 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__A2 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__I (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A2 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__A2 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__B1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__A1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__B1 (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A3 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__B1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__B2 (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__I (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__I (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__I (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__I (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__B (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A2 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__C (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__B (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__B2 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__I (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__I (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__I (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__B (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__B (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__B (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__B (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A2 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__A1 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__C (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__C (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__I (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__A1 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__A1 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A2 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__I (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A2 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A2 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__C (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__A1 (.I(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A1 (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A1 (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__A1 (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__I (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__B (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__B (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__A1 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A1 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A2 (.I(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__A2 (.I(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__A2 (.I(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__A2 (.I(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__B1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A2 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A2 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__B1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A1 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__B1 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__A2 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A2 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__A2 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__B1 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__B1 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__B1 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__B1 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__B1 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A1 (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__B (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11227__A1 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__B2 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__I (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__A1 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__I (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__B2 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__I (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A2 (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A1 (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__B1 (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__B (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__B2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__C1 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__C (.I(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__A1 (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A1 (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__I (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__A2 (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11594__I (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11581__A1 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A1 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A3 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__B (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__A2 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A2 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__C (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A1 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A2 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A2 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__I (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11588__A3 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__A3 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__B (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__B (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__B (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__B (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__I (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__A2 (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A2 (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__A2 (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__A2 (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__I (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__I (.I(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A2 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A2 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A2 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__A2 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__B2 (.I(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__B1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__B2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__B2 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__A2 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__A2 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A2 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__A2 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__B2 (.I(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A1 (.I(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A1 (.I(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__A1 (.I(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__A1 (.I(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__B2 (.I(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__B2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A2 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A2 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A2 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A2 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A1 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__A1 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A1 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A1 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__A2 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A2 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A2 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A2 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__B2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__B1 (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A2 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A2 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A2 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A2 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__B2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A2 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A2 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A2 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__A2 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__A1 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A1 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A1 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A1 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__B (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__B (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__B (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__I (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A2 (.I(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__A2 (.I(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A2 (.I(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A2 (.I(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A2 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__A2 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A2 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A2 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A1 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A1 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A1 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A1 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A2 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A2 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A2 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A2 (.I(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__A1 (.I(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A1 (.I(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__A1 (.I(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__A1 (.I(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A1 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__A1 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A1 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A1 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A1 (.I(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A1 (.I(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A1 (.I(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A1 (.I(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A1 (.I(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A1 (.I(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A1 (.I(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A1 (.I(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08825__A3 (.I(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__A3 (.I(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A2 (.I(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A2 (.I(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A2 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A2 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__I (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__I (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__I (.I(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__I (.I(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__I (.I(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__B (.I(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A2 (.I(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__I (.I(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__I (.I(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__I (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__C (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__I (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__I (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A3 (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__I (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__I (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__I (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__I (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A3 (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A4 (.I(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__I (.I(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A4 (.I(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A2 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A2 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A2 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A2 (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__C (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__I (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__I (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__I (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__B (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__B (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__I (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__I (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__I (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__I (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__I (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__I (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__B (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__I (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__B (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__I (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__I (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__I (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A2 (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A2 (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__A1 (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A2 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A4 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A2 (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A2 (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A2 (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A2 (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__I (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A2 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__I (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__I (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A3 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__I (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__I (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__B2 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__B2 (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__I (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__I (.I(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A2 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__A2 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A3 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A2 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__A2 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A2 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A2 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A2 (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A2 (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__B (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A2 (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__I (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__B (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__B (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A2 (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__B (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A1 (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A2 (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__C (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__C (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__S (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A1 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A1 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__B1 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__B1 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__B1 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__B1 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__B2 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__B (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A1 (.I(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A1 (.I(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A2 (.I(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A1 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__A1 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__A1 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A1 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A1 (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__A1 (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__A1 (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A1 (.I(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__A1 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A1 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A1 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__A1 (.I(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A1 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A1 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A2 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__B2 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__B2 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A2 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__A2 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__I (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__A1 (.I(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A1 (.I(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A2 (.I(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__B2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__C (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__B1 (.I(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__A2 (.I(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__B1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A2 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A1 (.I(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A1 (.I(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__B1 (.I(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A2 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__I (.I(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__I (.I(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A2 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A2 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A2 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A2 (.I(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__B2 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__B1 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__A1 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09328__A1 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A1 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A1 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A1 (.I(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__A1 (.I(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__A1 (.I(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A1 (.I(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A1 (.I(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__I (.I(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__I (.I(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__I (.I(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__I (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__I (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A2 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A2 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__S (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__S (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A1 (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A1 (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__I1 (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__B (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A1 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A1 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__I1 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A1 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__I0 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__I (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__S (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__S (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__S (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11222__A1 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A1 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__I1 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A1 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__I0 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A1 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A1 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__I1 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A1 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__I0 (.I(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__I1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A2 (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A2 (.I(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__I (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A2 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A2 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A2 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A2 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A1 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A1 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A2 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A2 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__A1 (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A1 (.I(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A2 (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A2 (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__A2 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A2 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A3 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__B1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__B1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A2 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__B1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__A2 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__A2 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__A2 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A2 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__A2 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A2 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__A1 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A2 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__A2 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11439__A2 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__B1 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A1 (.I(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__A1 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A1 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__A2 (.I(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A2 (.I(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A2 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__B1 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A3 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__A2 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11445__A2 (.I(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__B1 (.I(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__A1 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A1 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A1 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__A2 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A2 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A2 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__I (.I(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A2 (.I(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__B1 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09271__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__A3 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__I (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__A2 (.I(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__B1 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A1 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A1 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A2 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A2 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__A3 (.I(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__A2 (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A2 (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A1 (.I(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__B (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__A2 (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A2 (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__B (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__B (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__B (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__I (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09291__I (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__I (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__A2 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A2 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A2 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A2 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A2 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A2 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__A2 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A2 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A2 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A2 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A2 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__A2 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11416__A1 (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A1 (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A1 (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A1 (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__I (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__I (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__A2 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A2 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A2 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A2 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09328__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__B2 (.I(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__B1 (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__A1 (.I(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A1 (.I(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A1 (.I(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A1 (.I(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__B (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__B (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__B (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__I (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__I (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__I (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__A1 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A1 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__A1 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A1 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A1 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A1 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A1 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__A1 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__A1 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A1 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A1 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A1 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__A2 (.I(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A2 (.I(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A2 (.I(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A2 (.I(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A1 (.I(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A1 (.I(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A1 (.I(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A1 (.I(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__A1 (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A1 (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A1 (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__A1 (.I(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__B (.I(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__B (.I(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__B (.I(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__I (.I(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A2 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__A2 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__A2 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A2 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__I (.I(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__I (.I(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A2 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__A2 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__A2 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__A2 (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A2 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A2 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A2 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A2 (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__B2 (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__B1 (.I(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__A2 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__A2 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A2 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A2 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A2 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__A2 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A2 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A2 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__A2 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__B (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A1 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A2 (.I(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__S (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__I (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__I (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__S (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__S (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__S (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__S (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__A1 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A1 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A1 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__I1 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__B (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__B (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__B (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__I (.I(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__I (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__I (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A2 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A2 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A2 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A2 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__B2 (.I(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__B1 (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__A2 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A2 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A2 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A2 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__B (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__B (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__B (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__B (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A2 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A2 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A2 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A2 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A1 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A3 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__A3 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__A2 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__I (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__A2 (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__A1 (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__A1 (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A1 (.I(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__B (.I(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A2 (.I(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A1 (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__C (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__B (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__I (.I(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11588__A1 (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A1 (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A1 (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__B (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A3 (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A2 (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A1 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A1 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__B (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A1 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__A1 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A2 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A1 (.I(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__B (.I(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A3 (.I(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__B1 (.I(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A1 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__A2 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A3 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A2 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A3 (.I(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__B2 (.I(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__B1 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__B1 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__I (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__I (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A3 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__A1 (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__C (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__A1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__A1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__I (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__C (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__C (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A2 (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__B (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__C (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10681__I (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__I (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__I (.I(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__I (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__I (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A1 (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__A1 (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__B (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__B2 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__I (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__B2 (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__B2 (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__B2 (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A3 (.I(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A4 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A4 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A4 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__I1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__A2 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__B (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A2 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__A1 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__B (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A3 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A3 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__B1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__B1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A4 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__S (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__A1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__A3 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A1 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A3 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A1 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A1 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A1 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__A1 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__B (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__A2 (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A2 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__I (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__B (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A1 (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__C (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A4 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A3 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A3 (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A4 (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A2 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A4 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A2 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__A1 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A3 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A3 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A1 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A3 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__C (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A2 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__C (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A1 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__I (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A2 (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A1 (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A2 (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__A1 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A2 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A3 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__A2 (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A4 (.I(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__I (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__I (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__I (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__I (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__I (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__I (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__A1 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A1 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A1 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A1 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__A2 (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__A1 (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A1 (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__I (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__A1 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__A1 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__B (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A1 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__I (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A2 (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__I (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__I (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A1 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__A1 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__A1 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A1 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__B (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__B (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__I (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__B (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__B (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__C (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__B2 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A1 (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__A2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__A2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__I (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__I (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__A2 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A1 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__A1 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A2 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__B (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__C (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A1 (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A1 (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__B (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A2 (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__B (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__I (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__I (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__A2 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__B1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__B1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__B1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__A3 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A2 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__I (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__I (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__B (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__I (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__I (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__B1 (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__A1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__C (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__I (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__I (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__I (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A1 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__I (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__I (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A2 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A2 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A2 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__B (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__B (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__C (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__B (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__B2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__B2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__C (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__B (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__B (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A2 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__I (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__I (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__A3 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__B (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__I (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A1 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__A1 (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__B2 (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__B (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__B2 (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__B2 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__A1 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__B2 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__B1 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__C (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A1 (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__C (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__A1 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__I (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__B (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__B (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__I (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__C (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__C (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__C (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A1 (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11507__B (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__I (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__I (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__I (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__B2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11483__B (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__C (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__B (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__C (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__C (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__B (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__I (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__B1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__B2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__C (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__C (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__C (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__C (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__C (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__A2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A1 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__A1 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__C (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A1 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__A1 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A2 (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__A1 (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__B (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A1 (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A1 (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__A1 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__A1 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__B (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A1 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__A1 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09642__A1 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A1 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__I (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__A1 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__A1 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__A1 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A1 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A1 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__A2 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A2 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__A2 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A2 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__B2 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__A1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__B2 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__C (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__C (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__B (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__C (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A1 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11234__A1 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__A2 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A2 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A2 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__A1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__C (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09655__A1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__B2 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__A1 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__A1 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A2 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A2 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__A2 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A2 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__A2 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__C (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A2 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__B2 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__B2 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__B2 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__B2 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__C (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__C (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__C (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__B (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A1 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__C2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A1 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A1 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__A1 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A2 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__A2 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A2 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__B1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__A1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__A2 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A2 (.I(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A2 (.I(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__A1 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__B (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A2 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__I (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A2 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__A2 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__A2 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__B1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A3 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A2 (.I(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A2 (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__B1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__B1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11291__C (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__C (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__C (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__C (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A1 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__A2 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A2 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__A2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A1 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__I (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A1 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A2 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__A2 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A2 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__A2 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__I (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A2 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A2 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__A2 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__A2 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__A2 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__A2 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A1 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__B2 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__I (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__A2 (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A1 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__A1 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__A1 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__I (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A2 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A1 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A2 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__I (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__B2 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A2 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__I (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A3 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__B (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__C (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__B (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__C (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__A1 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__B2 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__A1 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A1 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__B (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A2 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__I (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__A2 (.I(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A1 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A2 (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A2 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A2 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__B1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__B1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__B1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__A1 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__C (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__B2 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__A1 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__A2 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__A2 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A1 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A1 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__A1 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__A2 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__C (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__C (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__C (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A1 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__A1 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A1 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A1 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__A2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A2 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__A1 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__A1 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__I (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__C (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A1 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__A1 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__C2 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__A1 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__A2 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A1 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A1 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__I (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A1 (.I(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A1 (.I(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__A2 (.I(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__B2 (.I(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__A2 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__A2 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A2 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A2 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A3 (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__B2 (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__B (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__B2 (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__A1 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11599__A1 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A1 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__B (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11139__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A2 (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__A2 (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__A2 (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A2 (.I(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__A1 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__A1 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__B2 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A1 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A1 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__A1 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__A1 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A1 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A2 (.I(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__A1 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A1 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__A1 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__I (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__I (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__B (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__A2 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__B2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__B2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__B2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A1 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__B1 (.I(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A2 (.I(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A2 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A2 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A1 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A1 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__B (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__B1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A1 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__C (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__C (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__B2 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A2 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10683__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A2 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A2 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__A1 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__B2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__C (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__A2 (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__A1 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__A1 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A1 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A1 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__B2 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__B2 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A1 (.I(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__A1 (.I(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A1 (.I(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__A1 (.I(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__B (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__A2 (.I(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A1 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__B2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A1 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A1 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__A2 (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__A2 (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A1 (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__B1 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__B (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__B (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A2 (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11584__C (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__C (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__C (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__B (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A1 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__A1 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__A1 (.I(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A2 (.I(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__A1 (.I(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__I (.I(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A2 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__I (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A1 (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__A1 (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A1 (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A1 (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A2 (.I(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A2 (.I(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__C (.I(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__B (.I(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__A2 (.I(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__A1 (.I(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__B2 (.I(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__A1 (.I(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__A1 (.I(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A2 (.I(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__A2 (.I(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__A1 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__A2 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__A2 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__A2 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A2 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__A2 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A2 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__A2 (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__A2 (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A1 (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A1 (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__B (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__A2 (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__A2 (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A2 (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__B (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__B (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__C (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__C (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__C (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A1 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__A1 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__B2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__A2 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A2 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__A2 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__B1 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__A1 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__A1 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__A1 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A1 (.I(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A2 (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__A1 (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A2 (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A1 (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A3 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__A2 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A3 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A2 (.I(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A2 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A2 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A3 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A2 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A3 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__A2 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__A1 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__A1 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__A1 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__B2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A2 (.I(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__A1 (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__B2 (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A1 (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A1 (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A2 (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__B1 (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__A1 (.I(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A2 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A2 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__A1 (.I(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A1 (.I(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A1 (.I(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__I (.I(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__A1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__A1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__I1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__B1 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11575__A1 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A1 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__B2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__B2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__A1 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__A1 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__A1 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A1 (.I(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__I (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A2 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A1 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A1 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__B2 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__A1 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__B (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__B (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__A1 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A1 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__A1 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A1 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__A1 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__A1 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__I (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__A1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__A1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__A2 (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A1 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__A1 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A1 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__B1 (.I(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__B1 (.I(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__A1 (.I(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__A1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__A1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__B1 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__B (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__C (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A1 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__A1 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A1 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__B2 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__A2 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A2 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__A2 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A1 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A1 (.I(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A1 (.I(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__A2 (.I(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__B (.I(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__A2 (.I(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A2 (.I(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__B2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__B1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__I (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__A1 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A1 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__A1 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__B2 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__A2 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A2 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A2 (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__A1 (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__A1 (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A1 (.I(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__A1 (.I(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__A1 (.I(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__A1 (.I(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__B2 (.I(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__A2 (.I(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A2 (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__B1 (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A2 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A2 (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A2 (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11548__B2 (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__B2 (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__C (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__B (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__B (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__B (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__B (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__B (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__A1 (.I(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A3 (.I(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__B (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__A2 (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A1 (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A3 (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__A2 (.I(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A2 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A3 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A2 (.I(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__A4 (.I(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__C (.I(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__A2 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__A2 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__A1 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__C (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__A1 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__I (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__B (.I(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A2 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__A1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__I (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__A1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__I (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__B (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__I (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__B2 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__I (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__A1 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__C (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__C (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A2 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__C (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__B (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__A2 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A1 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A4 (.I(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A2 (.I(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__A3 (.I(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__I (.I(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__A2 (.I(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__B1 (.I(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__B (.I(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__B (.I(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__A3 (.I(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A2 (.I(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A3 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__B (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A4 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__C (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A1 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A4 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__A2 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A4 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__A3 (.I(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A4 (.I(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__B1 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__B (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__I (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__C (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__I (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__C (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__B2 (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__C (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__B (.I(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__A2 (.I(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__B (.I(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__B (.I(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__I (.I(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__A1 (.I(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A2 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__A3 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__I (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__A1 (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__I (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__A1 (.I(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__B (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__A3 (.I(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__I (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__I (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__S (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__I (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__I (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__S (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A2 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A2 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A2 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__A2 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10915__A1 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__A1 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__A1 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A1 (.I(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A2 (.I(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__A2 (.I(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__A2 (.I(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A2 (.I(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__A2 (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__A1 (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A2 (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A1 (.I(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__B (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__A1 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__A1 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__A1 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__A1 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__A1 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__A2 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A1 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11620__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A1 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__I0 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A1 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A1 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A1 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__I1 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__I (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__I (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__I (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__I (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__C (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__C (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__C (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__C (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A3 (.I(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A2 (.I(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__A1 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A1 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A1 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A1 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A2 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__B (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__A2 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__B (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__A2 (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A1 (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A2 (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__I0 (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__C (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__C (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A1 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__I (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__C (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__C (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__C (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__A1 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__A2 (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__I (.I(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__I (.I(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__S (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A2 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__A2 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__S (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__I (.I(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__S (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__S (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__S (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__I (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__A1 (.I(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__A1 (.I(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__I (.I(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A2 (.I(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11617__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11544__B1 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11617__B (.I(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A2 (.I(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__A1 (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__A1 (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__C (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A2 (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A2 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__B (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A2 (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__A1 (.I(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__A1 (.I(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__A1 (.I(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__A2 (.I(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11613__A2 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__A2 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11613__B (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__A2 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11627__A2 (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__A2 (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__B (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11628__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11607__A2 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__I0 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__A2 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__I0 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A1 (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__A1 (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__A1 (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A1 (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A2 (.I(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__C (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__I (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__I (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A2 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__B1 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__A2 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A2 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__B1 (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__B1 (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__C (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__C (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__A1 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__A1 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__A1 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A2 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11588__A2 (.I(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__A1 (.I(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11528__A1 (.I(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A1 (.I(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11504__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__I (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__B2 (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__B (.I(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10867__I (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A2 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A1 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__I (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__C (.I(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A2 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__I (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__I (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__I (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__I (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__I (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__I (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__I (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A2 (.I(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11549__B (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11539__B (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__B (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__B (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__A2 (.I(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__C (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__C (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__C (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__C (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A2 (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A2 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A2 (.I(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A3 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A3 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__I (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__A2 (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A4 (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__I (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__I (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__I (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__C (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__I (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__B (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__I (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__A2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__A2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__A1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__A1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__I (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__B2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__B2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__I (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__I (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A1 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__I (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A1 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A1 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__A2 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__A2 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__B1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__B1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__A1 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__A1 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__A2 (.I(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__A2 (.I(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__B2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11507__A2 (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__C (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__C (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A1 (.I(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__S (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__A2 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__B2 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__B (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__B (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__I (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__A2 (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A2 (.I(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A3 (.I(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A2 (.I(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A2 (.I(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__A2 (.I(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__I (.I(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__A2 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__A2 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A2 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__A1 (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A1 (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10605__A1 (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A1 (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__A1 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A2 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__B (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__A2 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__I (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__A2 (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__A2 (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__A2 (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__A2 (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__A1 (.I(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__C (.I(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__B (.I(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__B (.I(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__A2 (.I(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A1 (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__A1 (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__A1 (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__A1 (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A2 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__A2 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__A1 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__I (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__I (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__I (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__A1 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__A1 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__A1 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A1 (.I(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__A2 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A2 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__A2 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__A1 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A1 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__C (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A1 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__C (.I(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__C (.I(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10607__C (.I(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__C (.I(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__B (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__S (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__I (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__I (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A1 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__A1 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A1 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__A1 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A1 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__A1 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__B (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A1 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__A2 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__A2 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__A4 (.I(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__B1 (.I(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__A2 (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__I (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A2 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__I (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A3 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A2 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__A2 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__A2 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__A2 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__B (.I(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__C (.I(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__C (.I(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__C (.I(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__C (.I(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__C (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__C (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__C (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__C (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__A2 (.I(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__A2 (.I(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__A1 (.I(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__A2 (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A2 (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__I (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__A2 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__A2 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A2 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__I (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__C (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A1 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__I (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11620__A1 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__A1 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__A1 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A1 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__A4 (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__A2 (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__B1 (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__A1 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A1 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__A1 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__A1 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A2 (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__B (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A1 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A1 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A1 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__A1 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A1 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__B (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__B1 (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__B (.I(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A2 (.I(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__A2 (.I(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__B1 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__B1 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__B1 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__A3 (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__A2 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11597__A2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__A2 (.I(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__B (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__A2 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A2 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10607__A2 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__A2 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__A2 (.I(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__A2 (.I(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A2 (.I(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__A2 (.I(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__A2 (.I(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A1 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A1 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__A1 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__A1 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10605__A4 (.I(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__A1 (.I(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__A2 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__A1 (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__A1 (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__B (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__C (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__B (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__A4 (.I(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10629__B (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__B1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__A2 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__A2 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__B1 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__C (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__C (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__C (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__C (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__A2 (.I(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__A2 (.I(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__A2 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__A2 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__A2 (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__I (.I(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__A2 (.I(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__A2 (.I(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__C (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A1 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10861__A1 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__C (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__B (.I(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A2 (.I(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__A2 (.I(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A4 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__A2 (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__B (.I(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__A1 (.I(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A2 (.I(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__B (.I(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__B (.I(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__B2 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__B2 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__B (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__C (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__A4 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A2 (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__B (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__A2 (.I(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__A2 (.I(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__B1 (.I(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__A2 (.I(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A2 (.I(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A2 (.I(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__A2 (.I(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__I (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__I (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__B2 (.I(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__A2 (.I(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__A2 (.I(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__A2 (.I(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__B2 (.I(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A1 (.I(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__A1 (.I(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__A1 (.I(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__C (.I(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__B (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A1 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__B (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A1 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A1 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__A2 (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A2 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__A2 (.I(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A1 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__A1 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A1 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A1 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__A1 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__B (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__A4 (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A2 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__B (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__C (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__C (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__C (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__A3 (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__A3 (.I(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11586__A2 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A2 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__B1 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A2 (.I(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__I (.I(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10737__I (.I(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__B2 (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A2 (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__B1 (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A2 (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__I1 (.I(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A2 (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A2 (.I(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__A2 (.I(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__A1 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A2 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__A4 (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__A2 (.I(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__A1 (.I(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A1 (.I(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A1 (.I(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__A1 (.I(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__A2 (.I(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__I (.I(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__I (.I(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__B2 (.I(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__A2 (.I(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__A2 (.I(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A2 (.I(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A1 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__A1 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A1 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__A1 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A1 (.I(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__B (.I(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__A2 (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__A2 (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__C (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__C (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__C (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__C (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__A1 (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A1 (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__B (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__B (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A2 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__C (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__B (.I(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__C (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__C (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__C (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__C (.I(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A2 (.I(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__B (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A3 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__C (.I(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__C (.I(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__C (.I(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__C (.I(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10809__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A2 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A2 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A2 (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__A2 (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A2 (.I(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__I (.I(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A2 (.I(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__A2 (.I(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A4 (.I(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__A2 (.I(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__A3 (.I(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__A2 (.I(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A2 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__B2 (.I(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A2 (.I(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__A2 (.I(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A2 (.I(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__A1 (.I(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__A2 (.I(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__A2 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__I (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__I (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__B2 (.I(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__A2 (.I(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__B1 (.I(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__A2 (.I(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__A1 (.I(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__B (.I(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__A1 (.I(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__A1 (.I(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__A3 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__A2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__A1 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A2 (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A2 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__A2 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__A3 (.I(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__A2 (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__B (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__B2 (.I(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__A2 (.I(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__A2 (.I(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A2 (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__B1 (.I(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A2 (.I(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__A2 (.I(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__A2 (.I(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__A2 (.I(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__C (.I(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A2 (.I(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__I (.I(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__A2 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__B2 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A1 (.I(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__A1 (.I(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A1 (.I(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__B2 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A2 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__A2 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A2 (.I(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A2 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A2 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__B1 (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A2 (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__A2 (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A3 (.I(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__B (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__B2 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A1 (.I(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A1 (.I(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A1 (.I(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A1 (.I(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__B2 (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A2 (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A2 (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A2 (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A2 (.I(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A2 (.I(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__A2 (.I(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A2 (.I(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__A1 (.I(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__B1 (.I(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A2 (.I(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A2 (.I(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A2 (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A2 (.I(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__C (.I(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__A2 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A2 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__B1 (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__B2 (.I(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__B1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A2 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__B1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__I (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A2 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__A3 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A2 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__A2 (.I(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A2 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A2 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11587__C (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__C (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__C (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__C (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__A2 (.I(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__I (.I(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__A2 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__A2 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__A2 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__A2 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A2 (.I(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__A2 (.I(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__B (.I(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__B1 (.I(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__B1 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__A1 (.I(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__I (.I(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__I (.I(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A3 (.I(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A4 (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11553__A1 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__A4 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A2 (.I(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__B (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A3 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A2 (.I(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__A1 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A3 (.I(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__I (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__I (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__I (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__I (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A1 (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A1 (.I(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A1 (.I(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__A1 (.I(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A1 (.I(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__A4 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__A2 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__A2 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A2 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__A2 (.I(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__B (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__A1 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A1 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__A2 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__C (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__C (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__A2 (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__A2 (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__C (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__A1 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__A1 (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__I (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__B (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__A1 (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__B (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__A1 (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__B1 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__B1 (.I(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__B1 (.I(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__B1 (.I(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__B1 (.I(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__B1 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__B1 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__B1 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__B1 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__I (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__I (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__C (.I(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__I (.I(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__I (.I(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__I (.I(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__A1 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A1 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A1 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__C (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11543__A2 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A2 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__A2 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__A2 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__B1 (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__B1 (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__B1 (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__B1 (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11075__I (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__I (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11510__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__I (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__I (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__C (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__A2 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A2 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__A2 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A2 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A2 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__B1 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__B1 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__B1 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__B1 (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__C (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__C (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__C (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__C (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__A2 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__A1 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__A1 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A1 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A2 (.I(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__B1 (.I(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__B1 (.I(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A2 (.I(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__C2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A2 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__A2 (.I(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11613__C (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__A1 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__C (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__C (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__A3 (.I(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__A2 (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A2 (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A1 (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A2 (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A2 (.I(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11533__B (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__B (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__B (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__C (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__A2 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__B1 (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__A2 (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__B1 (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__B1 (.I(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__A2 (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A2 (.I(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__A2 (.I(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A2 (.I(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A2 (.I(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__A2 (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A2 (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A2 (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A2 (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__C (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__C (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__C (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__I (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A1 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A1 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__A1 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11121__A1 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__A1 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11597__A1 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__B (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__A1 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A1 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__A1 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__B (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__B (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__A1 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__B1 (.I(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__C1 (.I(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__B1 (.I(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__B1 (.I(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A2 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__A2 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A2 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__A2 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__A2 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__A2 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__B1 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__B1 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__A2 (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__B2 (.I(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11139__A2 (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__A1 (.I(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A1 (.I(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__A1 (.I(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A1 (.I(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__B2 (.I(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11583__B (.I(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__C (.I(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__A2 (.I(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__C (.I(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A2 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__A1 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A1 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A1 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__B1 (.I(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__A1 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A1 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__B1 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__B1 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__A2 (.I(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__A2 (.I(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__B1 (.I(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A2 (.I(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A2 (.I(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__A2 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__A2 (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__B1 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11483__A1 (.I(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A1 (.I(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__A1 (.I(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__A1 (.I(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__B (.I(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__B (.I(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A1 (.I(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__A1 (.I(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__A2 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__A2 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A2 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A2 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__A2 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A2 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__A2 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A2 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__B1 (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__B1 (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__B1 (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__B1 (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A1 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__A2 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__C (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__C (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__C (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__C (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A2 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__B (.I(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__B1 (.I(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A2 (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__C2 (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A2 (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A2 (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A2 (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__A2 (.I(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__B1 (.I(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__B1 (.I(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__B1 (.I(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__A1 (.I(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__A1 (.I(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__C (.I(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__C (.I(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A2 (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__A2 (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A2 (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11208__A2 (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__B1 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__B1 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__B1 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11208__B1 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A2 (.I(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__B1 (.I(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__A1 (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__B1 (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__B1 (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__B1 (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__B1 (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A2 (.I(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11223__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__B (.I(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__B (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__A2 (.I(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A1 (.I(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A2 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__B1 (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__A1 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A2 (.I(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A2 (.I(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__A2 (.I(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A1 (.I(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__B (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A2 (.I(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__A1 (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__C (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A1 (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__B (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A2 (.I(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__B (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__A2 (.I(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__A3 (.I(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__A2 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A3 (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__A2 (.I(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__B (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__A2 (.I(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__B1 (.I(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__A2 (.I(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__B1 (.I(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__A2 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A2 (.I(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__A1 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__A1 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11586__A1 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A1 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__B1 (.I(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__B (.I(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__A4 (.I(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A2 (.I(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__A1 (.I(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__B1 (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__A3 (.I(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A2 (.I(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A3 (.I(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__A2 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__I (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__I (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__I (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__I (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__I (.I(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__A2 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A2 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__A2 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__A2 (.I(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__I (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__I (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__I (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__I (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__B (.I(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__B (.I(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__B (.I(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__C (.I(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__A2 (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__A2 (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A2 (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__A2 (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A2 (.I(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A2 (.I(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__A2 (.I(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__A2 (.I(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__B (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__B (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__B (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__B (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A2 (.I(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A2 (.I(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__A2 (.I(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__A2 (.I(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__B1 (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__A2 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__A2 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A2 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__A2 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A2 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__A2 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__A2 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__A2 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__A2 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11416__A2 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__A2 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__A2 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__A2 (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__A2 (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A2 (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__A2 (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__A2 (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__A2 (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__A2 (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__A2 (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__A2 (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__A2 (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__A3 (.I(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__B1 (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__B1 (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__B1 (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__B1 (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__A1 (.I(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__A1 (.I(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__A2 (.I(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__B1 (.I(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11467__A2 (.I(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__A2 (.I(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__A4 (.I(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__A2 (.I(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__B (.I(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11480__I (.I(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11548__A2 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__A1 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__A1 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11534__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__B (.I(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__A2 (.I(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A2 (.I(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__B1 (.I(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11527__I (.I(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__A2 (.I(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__A3 (.I(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11528__A3 (.I(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__A3 (.I(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__A2 (.I(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__A2 (.I(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__A2 (.I(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11528__A2 (.I(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11607__A1 (.I(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__B (.I(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11547__A2 (.I(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11537__A1 (.I(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11548__A1 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11544__A3 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__B1 (.I(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__A1 (.I(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__A1 (.I(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__B1 (.I(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__A2 (.I(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__I (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11591__A1 (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11563__A4 (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__B (.I(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__B (.I(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__A2 (.I(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__B (.I(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11575__A2 (.I(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__A2 (.I(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11587__A2 (.I(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11586__B (.I(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11585__A2 (.I(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11585__B (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11586__C (.I(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11591__A4 (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__B (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11592__A2 (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11596__A2 (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11617__A1 (.I(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11613__A1 (.I(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__A1 (.I(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__A1 (.I(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__A2 (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__A4 (.I(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__B (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__B (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11609__B2 (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__B (.I(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__C (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__I (.I(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A1 (.I(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A2 (.I(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05817__I (.I(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A2 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A1 (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__I (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05818__I (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11544__A1 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__A2 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A2 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__I (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A1 (.I(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A1 (.I(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__A1 (.I(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__I (.I(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__A1 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A1 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__B2 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__A1 (.I(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__A1 (.I(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__A2 (.I(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__A1 (.I(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__I (.I(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__A1 (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__I (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__A1 (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__I (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A1 (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__A1 (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__B (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__I (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__C (.I(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A2 (.I(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__I (.I(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__A1 (.I(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A2 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A2 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A1 (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05827__I (.I(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11502__I (.I(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__I (.I(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A1 (.I(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__A1 (.I(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__C2 (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__I (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__A1 (.I(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__S0 (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__S0 (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__A2 (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__I (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__I (.I(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__S0 (.I(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__S0 (.I(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__I (.I(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__I (.I(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__S0 (.I(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05843__A2 (.I(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__A2 (.I(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A1 (.I(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__I (.I(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05835__A1 (.I(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__I (.I(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__A1 (.I(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__I (.I(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05835__A2 (.I(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__A2 (.I(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__A2 (.I(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__I (.I(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__I (.I(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05847__A1 (.I(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05841__A1 (.I(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__I (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__A2 (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05847__A2 (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05840__I (.I(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A1 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__I (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A2 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__A3 (.I(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A1 (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A1 (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A1 (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05843__A1 (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__A1 (.I(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A1 (.I(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A1 (.I(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__A1 (.I(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A1 (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A1 (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__B1 (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__A1 (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__A2 (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05850__I (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__A1 (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A2 (.I(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__A2 (.I(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__B2 (.I(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__S (.I(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A1 (.I(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05984__A1 (.I(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__I (.I(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__A1 (.I(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__A1 (.I(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__A1 (.I(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__S0 (.I(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__S0 (.I(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__A2 (.I(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05852__A2 (.I(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__B2 (.I(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__B2 (.I(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__B2 (.I(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05862__A1 (.I(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__S (.I(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__S (.I(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__S (.I(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05857__I (.I(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__S1 (.I(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__S (.I(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__I (.I(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05859__I (.I(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__S1 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05892__S (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05867__S (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__I (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__I (.I(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__I (.I(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06480__A1 (.I(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__S1 (.I(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05862__A2 (.I(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__B2 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__B2 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__I (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__I (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__A1 (.I(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__I (.I(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__A1 (.I(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__A1 (.I(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A2 (.I(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A2 (.I(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__A2 (.I(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A1 (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A1 (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__A1 (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__I (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A1 (.I(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A1 (.I(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__I (.I(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A1 (.I(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A1 (.I(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__A2 (.I(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05890__A2 (.I(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__I (.I(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06480__A2 (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06192__I (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__A1 (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A2 (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06585__I (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__A1 (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A1 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A1 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A1 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05878__I (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A1 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A1 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__A1 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__I (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__A1 (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A1 (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__I (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__A1 (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__I (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__A2 (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__A2 (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__A2 (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__A1 (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__A1 (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__S1 (.I(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__S (.I(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__S1 (.I(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05883__S (.I(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A2 (.I(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A2 (.I(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__A2 (.I(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__B1 (.I(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__B2 (.I(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__C2 (.I(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__B2 (.I(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__B2 (.I(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__A1 (.I(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__A2 (.I(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__A2 (.I(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A1 (.I(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A1 (.I(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__A1 (.I(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__I (.I(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A1 (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__B2 (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07131__I (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05890__A1 (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A1 (.I(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__A1 (.I(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__A1 (.I(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__A1 (.I(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A2 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A2 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__A2 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__B1 (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__A1 (.I(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__A2 (.I(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__A2 (.I(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__I (.I(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05941__A2 (.I(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A4 (.I(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A1 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__A1 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A1 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__I (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__A1 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__A2 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__I (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__A1 (.I(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__S1 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__S (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__S1 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__S (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A2 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__A2 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__A2 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__B1 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__B1 (.I(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__C1 (.I(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__I (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__A1 (.I(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A1 (.I(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A1 (.I(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05906__I (.I(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__I (.I(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__A1 (.I(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__A1 (.I(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__A1 (.I(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__A2 (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__A2 (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__A2 (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__B1 (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__B1 (.I(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__C1 (.I(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A1 (.I(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A1 (.I(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07073__A1 (.I(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__I (.I(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__A1 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A1 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07112__A1 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__I (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__A1 (.I(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__I (.I(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__I (.I(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__A1 (.I(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__B1 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__B1 (.I(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__C1 (.I(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__I (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05956__A4 (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__A4 (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__I (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A4 (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__A1 (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__A2 (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__A3 (.I(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__I (.I(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__I (.I(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A1 (.I(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__A1 (.I(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A2 (.I(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__A1 (.I(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__A2 (.I(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__B2 (.I(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A1 (.I(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__A2 (.I(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05922__I (.I(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A1 (.I(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__A1 (.I(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__I (.I(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__A1 (.I(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__A2 (.I(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A1 (.I(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__A2 (.I(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__B1 (.I(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__B1 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__C1 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05970__I (.I(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__I (.I(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__A3 (.I(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A1 (.I(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__A1 (.I(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__I (.I(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__A1 (.I(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__A2 (.I(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__A2 (.I(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__A2 (.I(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__B1 (.I(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__B1 (.I(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__C1 (.I(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__I (.I(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__I (.I(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__A4 (.I(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__A2 (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__I1 (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05941__A3 (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A3 (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06136__A2 (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__A1 (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__A1 (.I(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__I (.I(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A1 (.I(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__A3 (.I(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A2 (.I(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A2 (.I(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A3 (.I(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A1 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A1 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__A1 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A1 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__A1 (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A1 (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A1 (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A2 (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07152__A1 (.I(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A1 (.I(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__I (.I(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__A1 (.I(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A1 (.I(_05806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__A2 (.I(_05806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A2 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__A2 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__A2 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__A1 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__A1 (.I(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A1 (.I(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A1 (.I(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__A1 (.I(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__I (.I(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__I (.I(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__I (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__I (.I(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__A2 (.I(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__A2 (.I(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A2 (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__I (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__A1 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__I (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__I (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__I (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05815__I (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__I (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A1 (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__I (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__I (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__I (.I(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__I (.I(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06175__A1 (.I(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__A1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__I (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__C (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__I1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__I1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__I (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__I1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__S0 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__A1 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05852__A1 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__I (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__A2 (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__A1 (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__A1 (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__I (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05934__A1 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__A1 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05825__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__A1 (.I(\as2650.ivec[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__I0 (.I(\as2650.ivec[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__A1 (.I(\as2650.ivec[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__I0 (.I(\as2650.ivec[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__A1 (.I(\as2650.ivec[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__I0 (.I(\as2650.ivec[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A1 (.I(\as2650.ivec[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__I0 (.I(\as2650.ivec[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__A1 (.I(\as2650.ivec[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__I0 (.I(\as2650.ivec[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__A1 (.I(\as2650.ivec[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__I0 (.I(\as2650.ivec[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A1 (.I(\as2650.ivec[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__I0 (.I(\as2650.ivec[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A1 (.I(\as2650.ivec[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A1 (.I(\as2650.ivec[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__A1 (.I(\as2650.last_intr ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A2 (.I(\as2650.last_intr ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__A2 (.I(\as2650.last_intr ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__I (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__I (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__I (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__I (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__I (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__I (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__I0 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__I1 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__I (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__I0 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__I1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__I (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__I0 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__I1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__I (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06917__I0 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__I1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__I (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__I0 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__I1 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__I (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__I0 (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__I1 (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__I (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__I0 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I1 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__I (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__I0 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__I1 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__A1 (.I(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__I0 (.I(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__A1 (.I(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__I0 (.I(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__A1 (.I(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__I0 (.I(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A1 (.I(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__I0 (.I(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__A1 (.I(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__I0 (.I(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A1 (.I(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I0 (.I(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A1 (.I(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__I0 (.I(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__B2 (.I(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05923__I0 (.I(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__B2 (.I(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__I0 (.I(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__B2 (.I(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__I0 (.I(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__B2 (.I(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__I0 (.I(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__I1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__I1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__I3 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__I1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__I3 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__I1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I3 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__I1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__I3 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__B2 (.I(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__I2 (.I(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__B2 (.I(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__I2 (.I(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__B2 (.I(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__I2 (.I(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__A1 (.I(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__I2 (.I(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__B2 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__B2 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A1 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__B2 (.I(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__B2 (.I(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A1 (.I(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__B2 (.I(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__B2 (.I(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A1 (.I(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__B2 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__B2 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A1 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__B2 (.I(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__B2 (.I(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__A1 (.I(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__B2 (.I(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__B2 (.I(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A1 (.I(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__A1 (.I(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__B2 (.I(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A1 (.I(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A1 (.I(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__B2 (.I(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A1 (.I(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A1 (.I(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__B2 (.I(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__A1 (.I(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__B2 (.I(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A1 (.I(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A1 (.I(\as2650.stack[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__C1 (.I(\as2650.stack[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A1 (.I(\as2650.stack[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__C1 (.I(\as2650.stack[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__A1 (.I(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__B2 (.I(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A1 (.I(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__C1 (.I(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__B2 (.I(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__A1 (.I(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A1 (.I(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__C1 (.I(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A1 (.I(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__A1 (.I(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__C1 (.I(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A1 (.I(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__C1 (.I(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__B2 (.I(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A1 (.I(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A1 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__B2 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A1 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__C1 (.I(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A1 (.I(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A1 (.I(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A1 (.I(\as2650.stack[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__A1 (.I(\as2650.stack[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__B2 (.I(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A1 (.I(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A1 (.I(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A1 (.I(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__C1 (.I(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__B2 (.I(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A1 (.I(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__A1 (.I(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__B2 (.I(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__A1 (.I(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__A1 (.I(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__B2 (.I(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A1 (.I(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A1 (.I(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__B2 (.I(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__A1 (.I(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A1 (.I(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__A1 (.I(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__A1 (.I(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A1 (.I(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__B2 (.I(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A1 (.I(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07766__A1 (.I(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__B2 (.I(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__C1 (.I(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A1 (.I(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A1 (.I(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__C1 (.I(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__B2 (.I(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__B2 (.I(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A1 (.I(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__A1 (.I(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__B2 (.I(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A1 (.I(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__B2 (.I(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A1 (.I(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__B2 (.I(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__B2 (.I(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__B2 (.I(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__A1 (.I(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__B2 (.I(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__B2 (.I(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A1 (.I(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__B2 (.I(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__B2 (.I(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A1 (.I(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__B2 (.I(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__B2 (.I(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A1 (.I(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__B2 (.I(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__B2 (.I(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__A1 (.I(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__B2 (.I(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__B2 (.I(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__A1 (.I(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11346__A1 (.I(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__B2 (.I(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A1 (.I(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A1 (.I(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__B2 (.I(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__A1 (.I(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__B2 (.I(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A1 (.I(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A1 (.I(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__A1 (.I(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__A1 (.I(\as2650.stack[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__B2 (.I(\as2650.stack[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__A1 (.I(\as2650.stack[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__B2 (.I(\as2650.stack[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__A1 (.I(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__A1 (.I(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A1 (.I(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A1 (.I(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__B2 (.I(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__A1 (.I(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__A1 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__A1 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__A1 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__A1 (.I(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A1 (.I(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__A1 (.I(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A1 (.I(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__A1 (.I(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__A1 (.I(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A1 (.I(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A1 (.I(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A1 (.I(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A1 (.I(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__B2 (.I(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__A1 (.I(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A1 (.I(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__B2 (.I(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A1 (.I(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__B2 (.I(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A1 (.I(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__B2 (.I(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A1 (.I(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A1 (.I(\as2650.stack[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A1 (.I(\as2650.stack[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__A1 (.I(\as2650.stack[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__A1 (.I(\as2650.stack[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A1 (.I(\as2650.stack[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A1 (.I(\as2650.stack[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A1 (.I(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__B2 (.I(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__A1 (.I(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A1 (.I(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__A1 (.I(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A1 (.I(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__A1 (.I(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__B2 (.I(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A1 (.I(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__A1 (.I(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__B2 (.I(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A1 (.I(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__A1 (.I(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__B2 (.I(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A1 (.I(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__A1 (.I(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__B2 (.I(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A1 (.I(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__C1 (.I(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A1 (.I(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A1 (.I(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A1 (.I(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A1 (.I(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__A1 (.I(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__A1 (.I(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__B2 (.I(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A1 (.I(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__A1 (.I(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__B2 (.I(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A1 (.I(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A1 (.I(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__B2 (.I(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__A1 (.I(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A1 (.I(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__B2 (.I(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__A1 (.I(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A1 (.I(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__B2 (.I(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__A1 (.I(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A1 (.I(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__B2 (.I(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A1 (.I(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__A1 (.I(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__A1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__A1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A1 (.I(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__C2 (.I(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__A1 (.I(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__C2 (.I(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A1 (.I(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__C2 (.I(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__A1 (.I(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__C2 (.I(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A1 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__A1 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A1 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A1 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__A1 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A1 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__A1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__B2 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__A1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__B2 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A1 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__B2 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__A1 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A1 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__A1 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A1 (.I(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__C2 (.I(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__A1 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__B2 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__A1 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__A1 (.I(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__A1 (.I(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A1 (.I(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A1 (.I(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__A1 (.I(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__A1 (.I(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A1 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__B2 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A1 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A1 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__A1 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A1 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__C1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__C1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__A1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A1 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__A1 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A1 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__A1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__C1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A1 (.I(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A1 (.I(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__A1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__B2 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A1 (.I(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A1 (.I(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A1 (.I(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A1 (.I(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A1 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A1 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A1 (.I(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A1 (.I(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__B2 (.I(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__A1 (.I(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A1 (.I(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__C2 (.I(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__A1 (.I(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__A1 (.I(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11208__B2 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__A1 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A1 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__B2 (.I(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__A1 (.I(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__A1 (.I(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__C2 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__B2 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__B2 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__C1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A1 (.I(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__A1 (.I(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A1 (.I(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__A1 (.I(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__B2 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__B2 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A1 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__A1 (.I(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__B2 (.I(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A1 (.I(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__B2 (.I(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A1 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__B2 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A1 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A1 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__B2 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A1 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__B2 (.I(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__B2 (.I(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A1 (.I(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__B2 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__B2 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__A1 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__A1 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__B2 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__A1 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__B2 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__A1 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__B2 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__B2 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__A1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__B2 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__A1 (.I(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__B2 (.I(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A1 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__A1 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A1 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A1 (.I(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__B2 (.I(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__A1 (.I(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__B2 (.I(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A1 (.I(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A1 (.I(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A1 (.I(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__A1 (.I(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A1 (.I(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A1 (.I(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__B2 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__B2 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A1 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A1 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__A1 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A1 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__A1 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__B2 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A1 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A1 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__B2 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A1 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__A1 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__B2 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A1 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__A1 (.I(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__A1 (.I(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A1 (.I(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__A1 (.I(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__A1 (.I(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__B2 (.I(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__A1 (.I(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A1 (.I(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A1 (.I(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A1 (.I(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A1 (.I(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A1 (.I(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__B2 (.I(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A1 (.I(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__B2 (.I(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A1 (.I(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__B2 (.I(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__A1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__C1 (.I(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__B2 (.I(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A1 (.I(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A1 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__A1 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__A1 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__A1 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__A1 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A1 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__C1 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__A1 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__A1 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__A1 (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A1 (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__B2 (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__B2 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A1 (.I(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__B2 (.I(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__A1 (.I(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__B2 (.I(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__B2 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__B2 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__B2 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__B2 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__A1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__A1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__B2 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A1 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A1 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__B2 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__A1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__B2 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A1 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A1 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__B2 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A1 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__A1 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A1 (.I(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__A1 (.I(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__B2 (.I(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__B2 (.I(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A1 (.I(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A1 (.I(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__B2 (.I(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A1 (.I(\as2650.stack[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__B2 (.I(\as2650.stack[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__B2 (.I(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__B2 (.I(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A1 (.I(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A1 (.I(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__B2 (.I(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A1 (.I(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__A1 (.I(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__B2 (.I(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__A1 (.I(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A1 (.I(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__B2 (.I(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A1 (.I(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__B2 (.I(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__B2 (.I(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A1 (.I(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__B2 (.I(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A1 (.I(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__B2 (.I(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__A1 (.I(\as2650.stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A1 (.I(\as2650.stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__B2 (.I(\as2650.stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A1 (.I(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__B2 (.I(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__A1 (.I(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A1 (.I(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A1 (.I(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__A1 (.I(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A1 (.I(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__A1 (.I(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__A1 (.I(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__A1 (.I(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__A1 (.I(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A1 (.I(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A1 (.I(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__A1 (.I(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__B2 (.I(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__A1 (.I(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A1 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__B2 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__A1 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A1 (.I(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A1 (.I(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__A1 (.I(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__A1 (.I(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__A1 (.I(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A1 (.I(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__A1 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A1 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A1 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06698__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output13_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__C2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output46_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A1 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output47_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output48_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11592__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__S (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__S (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output54_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A4 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output56_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A3 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__B (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A2 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output58_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output60_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output61_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output63_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07704__I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A2 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output66_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output67_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A1 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output69_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07332__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output71_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__A1 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output73_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07564__I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__B (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A2 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output74_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11629__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output75_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A3 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__A3 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output77_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A2 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__A2 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output79_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11093__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11622__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12131__I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output59_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A2 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output57_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output55_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__B2 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A3 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A2 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output53_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11648__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11804__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11809__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11721__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11810__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12041__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12040__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12048__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12038__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11961__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11957__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11955__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11962__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11990__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11995__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11991__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11633__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11635__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11862__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11832__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11831__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11834__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11835__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11858__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11645__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11869__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11866__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11828__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11641__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11637__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11631__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11634__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11639__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11938__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11871__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12023__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11870__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12022__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11971__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12027__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12026__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11636__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11972__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11970__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12025__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11951__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11950__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11974__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11922__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11945__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11854__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11845__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11946__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11943__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11942__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12032__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11940__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11941__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11933__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11936__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11934__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11932__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11925__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11926__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11930__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11931__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11929__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11898__CLK (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11899__CLK (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11918__CLK (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11903__CLK (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11904__CLK (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11905__CLK (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11900__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11902__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11914__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11915__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11901__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11989__CLK (.I(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11976__CLK (.I(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11975__CLK (.I(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11909__CLK (.I(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11986__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11985__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11987__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11984__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11983__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11757__CLK (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11758__CLK (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11765__CLK (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__CLK (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11763__CLK (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11760__CLK (.I(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11753__CLK (.I(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11752__CLK (.I(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11754__CLK (.I(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11755__CLK (.I(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11762__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11761__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11777__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11759__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11776__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11774__CLK (.I(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11788__CLK (.I(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11786__CLK (.I(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11787__CLK (.I(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11781__CLK (.I(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11783__CLK (.I(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__CLK (.I(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11725__CLK (.I(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11792__CLK (.I(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11794__CLK (.I(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11793__CLK (.I(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11782__CLK (.I(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11727__CLK (.I(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11729__CLK (.I(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11749__CLK (.I(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11751__CLK (.I(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11775__CLK (.I(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11769__CLK (.I(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__CLK (.I(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11767__CLK (.I(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11768__CLK (.I(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11916__CLK (.I(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11891__CLK (.I(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11764__CLK (.I(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__CLK (.I(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11897__CLK (.I(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11895__CLK (.I(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11896__CLK (.I(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__CLK (.I(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11877__CLK (.I(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11876__CLK (.I(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11824__CLK (.I(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12015__CLK (.I(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11825__CLK (.I(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11840__CLK (.I(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12017__CLK (.I(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12016__CLK (.I(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12018__CLK (.I(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11888__CLK (.I(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11889__CLK (.I(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__CLK (.I(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11841__CLK (.I(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12013__CLK (.I(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11827__CLK (.I(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11826__CLK (.I(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11736__CLK (.I(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11814__CLK (.I(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11737__CLK (.I(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11732__CLK (.I(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11735__CLK (.I(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11733__CLK (.I(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11812__CLK (.I(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__CLK (.I(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11816__CLK (.I(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11731__CLK (.I(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__CLK (.I(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11739__CLK (.I(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11724__CLK (.I(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11746__CLK (.I(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11750__CLK (.I(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11820__CLK (.I(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11704__CLK (.I(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11744__CLK (.I(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11743__CLK (.I(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11738__CLK (.I(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__CLK (.I(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__CLK (.I(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__CLK (.I(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11728__CLK (.I(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11741__CLK (.I(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11740__CLK (.I(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11742__CLK (.I(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11702__CLK (.I(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__CLK (.I(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12011__CLK (.I(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12006__CLK (.I(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12010__CLK (.I(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12009__CLK (.I(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12008__CLK (.I(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11797__CLK (.I(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11798__CLK (.I(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11695__CLK (.I(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12004__CLK (.I(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11800__CLK (.I(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11799__CLK (.I(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11665__CLK (.I(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11666__CLK (.I(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11664__CLK (.I(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__CLK (.I(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__CLK (.I(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11697__CLK (.I(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11795__CLK (.I(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11686__CLK (.I(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11657__CLK (.I(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11796__CLK (.I(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11658__CLK (.I(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__CLK (.I(clknet_leaf_131_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11673__CLK (.I(clknet_leaf_131_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__CLK (.I(clknet_leaf_131_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__CLK (.I(clknet_leaf_131_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11807__CLK (.I(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__CLK (.I(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11649__CLK (.I(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__CLK (.I(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11717__CLK (.I(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11650__CLK (.I(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11806__CLK (.I(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1_0_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0_0_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3_0_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2_0_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5_0_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4_0_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7_0_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6_0_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9_0_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8_0_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11_0_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10_0_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13_0_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12_0_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15_0_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14_0_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_132_wb_clk_i_I (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_131_wb_clk_i_I (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_130_wb_clk_i_I (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_129_wb_clk_i_I (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_128_wb_clk_i_I (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_126_wb_clk_i_I (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_wb_clk_i_I (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_wb_clk_i_I (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_122_wb_clk_i_I (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_wb_clk_i_I (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_135_wb_clk_i_I (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_134_wb_clk_i_I (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_133_wb_clk_i_I (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_wb_clk_i_I (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_wb_clk_i_I (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_wb_clk_i_I (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_wb_clk_i_I (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_wb_clk_i_I (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12012__CLK (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_wb_clk_i_I (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_wb_clk_i_I (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_wb_clk_i_I (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_wb_clk_i_I (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_wb_clk_i_I (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12007__CLK (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11789__CLK (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_wb_clk_i_I (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_wb_clk_i_I (.I(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_wb_clk_i_I (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_wb_clk_i_I (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_wb_clk_i_I (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_wb_clk_i_I (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_wb_clk_i_I (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_wb_clk_i_I (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_wb_clk_i_I (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_wb_clk_i_I (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_wb_clk_i_I (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_wb_clk_i_I (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11818__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11706__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12044__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12043__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12029__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11952__CLK (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11959__CLK (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11992__CLK (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11994__CLK (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11949__CLK (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11923__CLK (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11829__CLK (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11960__CLK (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_wb_clk_i_I (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_wb_clk_i_I (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_wb_clk_i_I (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_wb_clk_i_I (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_wb_clk_i_I (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11745__CLK (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_wb_clk_i_I (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_wb_clk_i_I (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_wb_clk_i_I (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_wb_clk_i_I (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_wb_clk_i_I (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_wb_clk_i_I (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_wb_clk_i_I (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_wb_clk_i_I (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_wb_clk_i_I (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_wb_clk_i_I (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_wb_clk_i_I (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_wb_clk_i_I (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12000__CLK (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_0_wb_clk_i_I (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_wb_clk_i_I (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_wb_clk_i_I (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11853__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11857__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11849__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11948__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_4_15_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__CLK (.I(clknet_4_15_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_4_15_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11999__CLK (.I(clknet_4_15_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_4_15_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_4_15_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12042__CLK (.I(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12001__CLK (.I(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1937 ();
 assign io_oeb[0] = net141;
 assign io_oeb[13] = net146;
 assign io_oeb[14] = net95;
 assign io_oeb[15] = net96;
 assign io_oeb[16] = net97;
 assign io_oeb[17] = net98;
 assign io_oeb[18] = net99;
 assign io_oeb[19] = net100;
 assign io_oeb[1] = net142;
 assign io_oeb[20] = net101;
 assign io_oeb[21] = net102;
 assign io_oeb[22] = net103;
 assign io_oeb[23] = net104;
 assign io_oeb[24] = net105;
 assign io_oeb[25] = net106;
 assign io_oeb[26] = net107;
 assign io_oeb[27] = net108;
 assign io_oeb[28] = net109;
 assign io_oeb[29] = net110;
 assign io_oeb[2] = net143;
 assign io_oeb[30] = net111;
 assign io_oeb[31] = net112;
 assign io_oeb[32] = net113;
 assign io_oeb[33] = net147;
 assign io_oeb[34] = net148;
 assign io_oeb[35] = net149;
 assign io_oeb[36] = net150;
 assign io_oeb[37] = net151;
 assign io_oeb[3] = net144;
 assign io_oeb[4] = net145;
 assign io_out[0] = net114;
 assign io_out[13] = net119;
 assign io_out[1] = net115;
 assign io_out[2] = net116;
 assign io_out[33] = net120;
 assign io_out[34] = net121;
 assign io_out[35] = net122;
 assign io_out[36] = net123;
 assign io_out[37] = net124;
 assign io_out[3] = net117;
 assign io_out[4] = net118;
 assign la_data_out[32] = net152;
 assign la_data_out[33] = net125;
 assign la_data_out[34] = net153;
 assign la_data_out[35] = net126;
 assign la_data_out[36] = net154;
 assign la_data_out[37] = net127;
 assign la_data_out[38] = net155;
 assign la_data_out[39] = net128;
 assign la_data_out[40] = net156;
 assign la_data_out[41] = net129;
 assign la_data_out[42] = net157;
 assign la_data_out[43] = net130;
 assign la_data_out[44] = net158;
 assign la_data_out[45] = net131;
 assign la_data_out[46] = net159;
 assign la_data_out[47] = net132;
 assign la_data_out[48] = net133;
 assign la_data_out[49] = net160;
 assign la_data_out[50] = net134;
 assign la_data_out[51] = net161;
 assign la_data_out[52] = net135;
 assign la_data_out[53] = net162;
 assign la_data_out[54] = net136;
 assign la_data_out[55] = net163;
 assign la_data_out[56] = net137;
 assign la_data_out[57] = net164;
 assign la_data_out[58] = net138;
 assign la_data_out[59] = net165;
 assign la_data_out[60] = net139;
 assign la_data_out[61] = net166;
 assign la_data_out[62] = net140;
 assign la_data_out[63] = net167;
endmodule

