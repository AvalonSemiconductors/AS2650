VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as2650
  CLASS BLOCK ;
  FOREIGN wrapped_as2650 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 700.000 ;
  PIN RAM_end_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 440.160 4.000 440.720 ;
    END
  END RAM_end_addr[0]
  PIN RAM_end_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 507.360 4.000 507.920 ;
    END
  END RAM_end_addr[10]
  PIN RAM_end_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 514.080 4.000 514.640 ;
    END
  END RAM_end_addr[11]
  PIN RAM_end_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 520.800 4.000 521.360 ;
    END
  END RAM_end_addr[12]
  PIN RAM_end_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 527.520 4.000 528.080 ;
    END
  END RAM_end_addr[13]
  PIN RAM_end_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 534.240 4.000 534.800 ;
    END
  END RAM_end_addr[14]
  PIN RAM_end_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 540.960 4.000 541.520 ;
    END
  END RAM_end_addr[15]
  PIN RAM_end_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 446.880 4.000 447.440 ;
    END
  END RAM_end_addr[1]
  PIN RAM_end_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 453.600 4.000 454.160 ;
    END
  END RAM_end_addr[2]
  PIN RAM_end_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 460.320 4.000 460.880 ;
    END
  END RAM_end_addr[3]
  PIN RAM_end_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 467.040 4.000 467.600 ;
    END
  END RAM_end_addr[4]
  PIN RAM_end_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 473.760 4.000 474.320 ;
    END
  END RAM_end_addr[5]
  PIN RAM_end_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 480.480 4.000 481.040 ;
    END
  END RAM_end_addr[6]
  PIN RAM_end_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 487.200 4.000 487.760 ;
    END
  END RAM_end_addr[7]
  PIN RAM_end_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 493.920 4.000 494.480 ;
    END
  END RAM_end_addr[8]
  PIN RAM_end_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 500.640 4.000 501.200 ;
    END
  END RAM_end_addr[9]
  PIN RAM_start_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 305.760 4.000 306.320 ;
    END
  END RAM_start_addr[0]
  PIN RAM_start_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 372.960 4.000 373.520 ;
    END
  END RAM_start_addr[10]
  PIN RAM_start_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 379.680 4.000 380.240 ;
    END
  END RAM_start_addr[11]
  PIN RAM_start_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.400 4.000 386.960 ;
    END
  END RAM_start_addr[12]
  PIN RAM_start_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 393.120 4.000 393.680 ;
    END
  END RAM_start_addr[13]
  PIN RAM_start_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 399.840 4.000 400.400 ;
    END
  END RAM_start_addr[14]
  PIN RAM_start_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 406.560 4.000 407.120 ;
    END
  END RAM_start_addr[15]
  PIN RAM_start_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 312.480 4.000 313.040 ;
    END
  END RAM_start_addr[1]
  PIN RAM_start_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.200 4.000 319.760 ;
    END
  END RAM_start_addr[2]
  PIN RAM_start_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 325.920 4.000 326.480 ;
    END
  END RAM_start_addr[3]
  PIN RAM_start_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 332.640 4.000 333.200 ;
    END
  END RAM_start_addr[4]
  PIN RAM_start_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 339.360 4.000 339.920 ;
    END
  END RAM_start_addr[5]
  PIN RAM_start_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 346.080 4.000 346.640 ;
    END
  END RAM_start_addr[6]
  PIN RAM_start_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.800 4.000 353.360 ;
    END
  END RAM_start_addr[7]
  PIN RAM_start_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 359.520 4.000 360.080 ;
    END
  END RAM_start_addr[8]
  PIN RAM_start_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 366.240 4.000 366.800 ;
    END
  END RAM_start_addr[9]
  PIN WEb_raw
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 946.400 696.000 946.960 700.000 ;
    END
  END WEb_raw
  PIN boot_rom_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 433.440 4.000 434.000 ;
    END
  END boot_rom_en
  PIN bus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 679.840 696.000 680.400 700.000 ;
    END
  END bus_addr[0]
  PIN bus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 696.000 699.440 700.000 ;
    END
  END bus_addr[1]
  PIN bus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 717.920 696.000 718.480 700.000 ;
    END
  END bus_addr[2]
  PIN bus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 736.960 696.000 737.520 700.000 ;
    END
  END bus_addr[3]
  PIN bus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 756.000 696.000 756.560 700.000 ;
    END
  END bus_addr[4]
  PIN bus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 775.040 696.000 775.600 700.000 ;
    END
  END bus_addr[5]
  PIN bus_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 660.800 696.000 661.360 700.000 ;
    END
  END bus_cyc
  PIN bus_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 696.000 509.040 700.000 ;
    END
  END bus_data_out[0]
  PIN bus_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 696.000 528.080 700.000 ;
    END
  END bus_data_out[1]
  PIN bus_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 546.560 696.000 547.120 700.000 ;
    END
  END bus_data_out[2]
  PIN bus_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 565.600 696.000 566.160 700.000 ;
    END
  END bus_data_out[3]
  PIN bus_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 696.000 585.200 700.000 ;
    END
  END bus_data_out[4]
  PIN bus_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 603.680 696.000 604.240 700.000 ;
    END
  END bus_data_out[5]
  PIN bus_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 622.720 696.000 623.280 700.000 ;
    END
  END bus_data_out[6]
  PIN bus_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 696.000 642.320 700.000 ;
    END
  END bus_data_out[7]
  PIN bus_in_gpios[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 514.080 1000.000 514.640 ;
    END
  END bus_in_gpios[0]
  PIN bus_in_gpios[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 521.920 1000.000 522.480 ;
    END
  END bus_in_gpios[1]
  PIN bus_in_gpios[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 529.760 1000.000 530.320 ;
    END
  END bus_in_gpios[2]
  PIN bus_in_gpios[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 537.600 1000.000 538.160 ;
    END
  END bus_in_gpios[3]
  PIN bus_in_gpios[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 545.440 1000.000 546.000 ;
    END
  END bus_in_gpios[4]
  PIN bus_in_gpios[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 553.280 1000.000 553.840 ;
    END
  END bus_in_gpios[5]
  PIN bus_in_gpios[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 561.120 1000.000 561.680 ;
    END
  END bus_in_gpios[6]
  PIN bus_in_gpios[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 568.960 1000.000 569.520 ;
    END
  END bus_in_gpios[7]
  PIN bus_in_serial_ports[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 794.080 696.000 794.640 700.000 ;
    END
  END bus_in_serial_ports[0]
  PIN bus_in_serial_ports[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 696.000 813.680 700.000 ;
    END
  END bus_in_serial_ports[1]
  PIN bus_in_serial_ports[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 832.160 696.000 832.720 700.000 ;
    END
  END bus_in_serial_ports[2]
  PIN bus_in_serial_ports[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 851.200 696.000 851.760 700.000 ;
    END
  END bus_in_serial_ports[3]
  PIN bus_in_serial_ports[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 696.000 870.800 700.000 ;
    END
  END bus_in_serial_ports[4]
  PIN bus_in_serial_ports[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 889.280 696.000 889.840 700.000 ;
    END
  END bus_in_serial_ports[5]
  PIN bus_in_serial_ports[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 908.320 696.000 908.880 700.000 ;
    END
  END bus_in_serial_ports[6]
  PIN bus_in_serial_ports[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 696.000 927.920 700.000 ;
    END
  END bus_in_serial_ports[7]
  PIN bus_in_timers[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 600.320 1000.000 600.880 ;
    END
  END bus_in_timers[0]
  PIN bus_in_timers[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 608.160 1000.000 608.720 ;
    END
  END bus_in_timers[1]
  PIN bus_in_timers[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 616.000 1000.000 616.560 ;
    END
  END bus_in_timers[2]
  PIN bus_in_timers[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 623.840 1000.000 624.400 ;
    END
  END bus_in_timers[3]
  PIN bus_in_timers[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 631.680 1000.000 632.240 ;
    END
  END bus_in_timers[4]
  PIN bus_in_timers[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 639.520 1000.000 640.080 ;
    END
  END bus_in_timers[5]
  PIN bus_in_timers[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 647.360 1000.000 647.920 ;
    END
  END bus_in_timers[6]
  PIN bus_in_timers[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 655.200 1000.000 655.760 ;
    END
  END bus_in_timers[7]
  PIN bus_we_gpios
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 506.240 1000.000 506.800 ;
    END
  END bus_we_gpios
  PIN bus_we_serial_ports
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 592.480 1000.000 593.040 ;
    END
  END bus_we_serial_ports
  PIN bus_we_timers
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 584.640 1000.000 585.200 ;
    END
  END bus_we_timers
  PIN cs_port[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 413.280 4.000 413.840 ;
    END
  END cs_port[0]
  PIN cs_port[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 420.000 4.000 420.560 ;
    END
  END cs_port[1]
  PIN cs_port[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 426.720 4.000 427.280 ;
    END
  END cs_port[2]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 696.000 14.000 700.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 696.000 204.400 700.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 696.000 223.440 700.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 696.000 242.480 700.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 696.000 261.520 700.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 696.000 280.560 700.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 696.000 299.600 700.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.080 696.000 318.640 700.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 696.000 337.680 700.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 696.000 356.720 700.000 ;
    END
  END io_in[18]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 696.000 33.040 700.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 696.000 52.080 700.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 696.000 71.120 700.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 696.000 90.160 700.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 696.000 109.200 700.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 696.000 128.240 700.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 696.000 147.280 700.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 696.000 166.320 700.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 696.000 185.360 700.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 4.000 178.640 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 245.280 4.000 245.840 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 4.000 252.560 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.720 4.000 259.280 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 265.440 4.000 266.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 272.160 4.000 272.720 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.880 4.000 279.440 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.600 4.000 286.160 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 292.320 4.000 292.880 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 299.040 4.000 299.600 ;
    END
  END io_oeb[18]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 4.000 192.080 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.240 4.000 198.800 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 4.000 205.520 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 4.000 212.240 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 4.000 218.960 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.120 4.000 225.680 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 231.840 4.000 232.400 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 4.000 239.120 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.400 4.000 50.960 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 171.360 4.000 171.920 ;
    END
  END io_out[18]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 4.000 57.680 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.840 4.000 64.400 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 4.000 71.120 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.280 4.000 77.840 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 4.000 84.560 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.440 4.000 98.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 482.720 1000.000 483.280 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 490.560 1000.000 491.120 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 498.400 1000.000 498.960 ;
    END
  END irq[2]
  PIN irqs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 696.000 375.760 700.000 ;
    END
  END irqs[0]
  PIN irqs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 394.240 696.000 394.800 700.000 ;
    END
  END irqs[1]
  PIN irqs[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 696.000 413.840 700.000 ;
    END
  END irqs[2]
  PIN irqs[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 696.000 432.880 700.000 ;
    END
  END irqs[3]
  PIN irqs[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 696.000 451.920 700.000 ;
    END
  END irqs[4]
  PIN irqs[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 696.000 470.960 700.000 ;
    END
  END irqs[5]
  PIN irqs[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 489.440 696.000 490.000 700.000 ;
    END
  END irqs[6]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 43.680 1000.000 44.240 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 122.080 1000.000 122.640 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 129.920 1000.000 130.480 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 137.760 1000.000 138.320 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 145.600 1000.000 146.160 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 153.440 1000.000 154.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 161.280 1000.000 161.840 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 169.120 1000.000 169.680 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 176.960 1000.000 177.520 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 184.800 1000.000 185.360 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 192.640 1000.000 193.200 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 51.520 1000.000 52.080 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 200.480 1000.000 201.040 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 208.320 1000.000 208.880 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 216.160 1000.000 216.720 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 224.000 1000.000 224.560 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 231.840 1000.000 232.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 239.680 1000.000 240.240 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 247.520 1000.000 248.080 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 255.360 1000.000 255.920 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 263.200 1000.000 263.760 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 271.040 1000.000 271.600 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 59.360 1000.000 59.920 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 278.880 1000.000 279.440 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 286.720 1000.000 287.280 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 294.560 1000.000 295.120 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 302.400 1000.000 302.960 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 310.240 1000.000 310.800 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 318.080 1000.000 318.640 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 325.920 1000.000 326.480 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 333.760 1000.000 334.320 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 341.600 1000.000 342.160 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 349.440 1000.000 350.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 67.200 1000.000 67.760 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 357.280 1000.000 357.840 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 365.120 1000.000 365.680 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 372.960 1000.000 373.520 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 380.800 1000.000 381.360 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 388.640 1000.000 389.200 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 396.480 1000.000 397.040 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 404.320 1000.000 404.880 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 412.160 1000.000 412.720 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 420.000 1000.000 420.560 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 427.840 1000.000 428.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 75.040 1000.000 75.600 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 435.680 1000.000 436.240 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 443.520 1000.000 444.080 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 451.360 1000.000 451.920 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 459.200 1000.000 459.760 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 467.040 1000.000 467.600 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 474.880 1000.000 475.440 ;
    END
  END la_data_out[55]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 82.880 1000.000 83.440 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 90.720 1000.000 91.280 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 98.560 1000.000 99.120 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 106.400 1000.000 106.960 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 114.240 1000.000 114.800 ;
    END
  END la_data_out[9]
  PIN le_hi_act
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 696.000 985.040 700.000 ;
    END
  END le_hi_act
  PIN le_lo_act
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 965.440 696.000 966.000 700.000 ;
    END
  END le_lo_act
  PIN reset_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 576.800 1000.000 577.360 ;
    END
  END reset_out
  PIN rom_bus_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 601.440 4.000 602.000 ;
    END
  END rom_bus_in[0]
  PIN rom_bus_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 608.160 4.000 608.720 ;
    END
  END rom_bus_in[1]
  PIN rom_bus_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 614.880 4.000 615.440 ;
    END
  END rom_bus_in[2]
  PIN rom_bus_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 621.600 4.000 622.160 ;
    END
  END rom_bus_in[3]
  PIN rom_bus_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 628.320 4.000 628.880 ;
    END
  END rom_bus_in[4]
  PIN rom_bus_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 635.040 4.000 635.600 ;
    END
  END rom_bus_in[5]
  PIN rom_bus_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 641.760 4.000 642.320 ;
    END
  END rom_bus_in[6]
  PIN rom_bus_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 648.480 4.000 649.040 ;
    END
  END rom_bus_in[7]
  PIN rom_bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 547.680 4.000 548.240 ;
    END
  END rom_bus_out[0]
  PIN rom_bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 554.400 4.000 554.960 ;
    END
  END rom_bus_out[1]
  PIN rom_bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 561.120 4.000 561.680 ;
    END
  END rom_bus_out[2]
  PIN rom_bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 567.840 4.000 568.400 ;
    END
  END rom_bus_out[3]
  PIN rom_bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.560 4.000 575.120 ;
    END
  END rom_bus_out[4]
  PIN rom_bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 581.280 4.000 581.840 ;
    END
  END rom_bus_out[5]
  PIN rom_bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 588.000 4.000 588.560 ;
    END
  END rom_bus_out[6]
  PIN rom_bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 594.720 4.000 595.280 ;
    END
  END rom_bus_out[7]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 682.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 682.380 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 0.000 65.520 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 0.000 370.160 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 0.000 397.040 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 0.000 423.920 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 0.000 450.800 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 0.000 477.680 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 0.000 504.560 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 0.000 531.440 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 0.000 558.320 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 0.000 585.200 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 0.000 612.080 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 0.000 638.960 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 0.000 665.840 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 0.000 692.720 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 0.000 719.600 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 0.000 746.480 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 0.000 773.360 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 0.000 800.240 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 826.560 0.000 827.120 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 853.440 0.000 854.000 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 880.320 0.000 880.880 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 0.000 907.760 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 934.080 0.000 934.640 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 0.000 182.000 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 0.000 208.880 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 0.000 235.760 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 0.000 262.640 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 0.000 289.520 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 0.000 316.400 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 0.000 343.280 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 0.000 110.320 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 0.000 379.120 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 405.440 0.000 406.000 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 0.000 432.880 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 0.000 459.760 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 486.080 0.000 486.640 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 512.960 0.000 513.520 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 0.000 540.400 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 566.720 0.000 567.280 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 593.600 0.000 594.160 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 620.480 0.000 621.040 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 0.000 137.200 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 647.360 0.000 647.920 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 674.240 0.000 674.800 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 701.120 0.000 701.680 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 728.000 0.000 728.560 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 754.880 0.000 755.440 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 781.760 0.000 782.320 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 808.640 0.000 809.200 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 835.520 0.000 836.080 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 0.000 862.960 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 889.280 0.000 889.840 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 0.000 164.080 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 916.160 0.000 916.720 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 943.040 0.000 943.600 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 0.000 190.960 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 0.000 217.840 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 0.000 244.720 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 0.000 271.600 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 0.000 298.480 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 0.000 325.360 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 0.000 352.240 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 0.000 119.280 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 0.000 388.080 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 0.000 414.960 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 0.000 441.840 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 468.160 0.000 468.720 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 495.040 0.000 495.600 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 521.920 0.000 522.480 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 0.000 549.360 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 0.000 576.240 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 602.560 0.000 603.120 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 629.440 0.000 630.000 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 0.000 146.160 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 656.320 0.000 656.880 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 683.200 0.000 683.760 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 710.080 0.000 710.640 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 736.960 0.000 737.520 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 763.840 0.000 764.400 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 790.720 0.000 791.280 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 817.600 0.000 818.160 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 844.480 0.000 845.040 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 871.360 0.000 871.920 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 898.240 0.000 898.800 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 0.000 173.040 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 925.120 0.000 925.680 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 952.000 0.000 952.560 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 0.000 199.920 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 0.000 253.680 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 0.000 280.560 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 0.000 307.440 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 0.000 334.320 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 0.000 361.200 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 0.000 83.440 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 0.000 92.400 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 992.880 682.380 ;
      LAYER Metal2 ;
        RECT 6.860 695.700 13.140 696.500 ;
        RECT 14.300 695.700 32.180 696.500 ;
        RECT 33.340 695.700 51.220 696.500 ;
        RECT 52.380 695.700 70.260 696.500 ;
        RECT 71.420 695.700 89.300 696.500 ;
        RECT 90.460 695.700 108.340 696.500 ;
        RECT 109.500 695.700 127.380 696.500 ;
        RECT 128.540 695.700 146.420 696.500 ;
        RECT 147.580 695.700 165.460 696.500 ;
        RECT 166.620 695.700 184.500 696.500 ;
        RECT 185.660 695.700 203.540 696.500 ;
        RECT 204.700 695.700 222.580 696.500 ;
        RECT 223.740 695.700 241.620 696.500 ;
        RECT 242.780 695.700 260.660 696.500 ;
        RECT 261.820 695.700 279.700 696.500 ;
        RECT 280.860 695.700 298.740 696.500 ;
        RECT 299.900 695.700 317.780 696.500 ;
        RECT 318.940 695.700 336.820 696.500 ;
        RECT 337.980 695.700 355.860 696.500 ;
        RECT 357.020 695.700 374.900 696.500 ;
        RECT 376.060 695.700 393.940 696.500 ;
        RECT 395.100 695.700 412.980 696.500 ;
        RECT 414.140 695.700 432.020 696.500 ;
        RECT 433.180 695.700 451.060 696.500 ;
        RECT 452.220 695.700 470.100 696.500 ;
        RECT 471.260 695.700 489.140 696.500 ;
        RECT 490.300 695.700 508.180 696.500 ;
        RECT 509.340 695.700 527.220 696.500 ;
        RECT 528.380 695.700 546.260 696.500 ;
        RECT 547.420 695.700 565.300 696.500 ;
        RECT 566.460 695.700 584.340 696.500 ;
        RECT 585.500 695.700 603.380 696.500 ;
        RECT 604.540 695.700 622.420 696.500 ;
        RECT 623.580 695.700 641.460 696.500 ;
        RECT 642.620 695.700 660.500 696.500 ;
        RECT 661.660 695.700 679.540 696.500 ;
        RECT 680.700 695.700 698.580 696.500 ;
        RECT 699.740 695.700 717.620 696.500 ;
        RECT 718.780 695.700 736.660 696.500 ;
        RECT 737.820 695.700 755.700 696.500 ;
        RECT 756.860 695.700 774.740 696.500 ;
        RECT 775.900 695.700 793.780 696.500 ;
        RECT 794.940 695.700 812.820 696.500 ;
        RECT 813.980 695.700 831.860 696.500 ;
        RECT 833.020 695.700 850.900 696.500 ;
        RECT 852.060 695.700 869.940 696.500 ;
        RECT 871.100 695.700 888.980 696.500 ;
        RECT 890.140 695.700 908.020 696.500 ;
        RECT 909.180 695.700 927.060 696.500 ;
        RECT 928.220 695.700 946.100 696.500 ;
        RECT 947.260 695.700 965.140 696.500 ;
        RECT 966.300 695.700 984.180 696.500 ;
        RECT 985.340 695.700 994.420 696.500 ;
        RECT 6.860 4.300 994.420 695.700 ;
        RECT 6.860 3.500 46.740 4.300 ;
        RECT 47.900 3.500 55.700 4.300 ;
        RECT 56.860 3.500 64.660 4.300 ;
        RECT 65.820 3.500 73.620 4.300 ;
        RECT 74.780 3.500 82.580 4.300 ;
        RECT 83.740 3.500 91.540 4.300 ;
        RECT 92.700 3.500 100.500 4.300 ;
        RECT 101.660 3.500 109.460 4.300 ;
        RECT 110.620 3.500 118.420 4.300 ;
        RECT 119.580 3.500 127.380 4.300 ;
        RECT 128.540 3.500 136.340 4.300 ;
        RECT 137.500 3.500 145.300 4.300 ;
        RECT 146.460 3.500 154.260 4.300 ;
        RECT 155.420 3.500 163.220 4.300 ;
        RECT 164.380 3.500 172.180 4.300 ;
        RECT 173.340 3.500 181.140 4.300 ;
        RECT 182.300 3.500 190.100 4.300 ;
        RECT 191.260 3.500 199.060 4.300 ;
        RECT 200.220 3.500 208.020 4.300 ;
        RECT 209.180 3.500 216.980 4.300 ;
        RECT 218.140 3.500 225.940 4.300 ;
        RECT 227.100 3.500 234.900 4.300 ;
        RECT 236.060 3.500 243.860 4.300 ;
        RECT 245.020 3.500 252.820 4.300 ;
        RECT 253.980 3.500 261.780 4.300 ;
        RECT 262.940 3.500 270.740 4.300 ;
        RECT 271.900 3.500 279.700 4.300 ;
        RECT 280.860 3.500 288.660 4.300 ;
        RECT 289.820 3.500 297.620 4.300 ;
        RECT 298.780 3.500 306.580 4.300 ;
        RECT 307.740 3.500 315.540 4.300 ;
        RECT 316.700 3.500 324.500 4.300 ;
        RECT 325.660 3.500 333.460 4.300 ;
        RECT 334.620 3.500 342.420 4.300 ;
        RECT 343.580 3.500 351.380 4.300 ;
        RECT 352.540 3.500 360.340 4.300 ;
        RECT 361.500 3.500 369.300 4.300 ;
        RECT 370.460 3.500 378.260 4.300 ;
        RECT 379.420 3.500 387.220 4.300 ;
        RECT 388.380 3.500 396.180 4.300 ;
        RECT 397.340 3.500 405.140 4.300 ;
        RECT 406.300 3.500 414.100 4.300 ;
        RECT 415.260 3.500 423.060 4.300 ;
        RECT 424.220 3.500 432.020 4.300 ;
        RECT 433.180 3.500 440.980 4.300 ;
        RECT 442.140 3.500 449.940 4.300 ;
        RECT 451.100 3.500 458.900 4.300 ;
        RECT 460.060 3.500 467.860 4.300 ;
        RECT 469.020 3.500 476.820 4.300 ;
        RECT 477.980 3.500 485.780 4.300 ;
        RECT 486.940 3.500 494.740 4.300 ;
        RECT 495.900 3.500 503.700 4.300 ;
        RECT 504.860 3.500 512.660 4.300 ;
        RECT 513.820 3.500 521.620 4.300 ;
        RECT 522.780 3.500 530.580 4.300 ;
        RECT 531.740 3.500 539.540 4.300 ;
        RECT 540.700 3.500 548.500 4.300 ;
        RECT 549.660 3.500 557.460 4.300 ;
        RECT 558.620 3.500 566.420 4.300 ;
        RECT 567.580 3.500 575.380 4.300 ;
        RECT 576.540 3.500 584.340 4.300 ;
        RECT 585.500 3.500 593.300 4.300 ;
        RECT 594.460 3.500 602.260 4.300 ;
        RECT 603.420 3.500 611.220 4.300 ;
        RECT 612.380 3.500 620.180 4.300 ;
        RECT 621.340 3.500 629.140 4.300 ;
        RECT 630.300 3.500 638.100 4.300 ;
        RECT 639.260 3.500 647.060 4.300 ;
        RECT 648.220 3.500 656.020 4.300 ;
        RECT 657.180 3.500 664.980 4.300 ;
        RECT 666.140 3.500 673.940 4.300 ;
        RECT 675.100 3.500 682.900 4.300 ;
        RECT 684.060 3.500 691.860 4.300 ;
        RECT 693.020 3.500 700.820 4.300 ;
        RECT 701.980 3.500 709.780 4.300 ;
        RECT 710.940 3.500 718.740 4.300 ;
        RECT 719.900 3.500 727.700 4.300 ;
        RECT 728.860 3.500 736.660 4.300 ;
        RECT 737.820 3.500 745.620 4.300 ;
        RECT 746.780 3.500 754.580 4.300 ;
        RECT 755.740 3.500 763.540 4.300 ;
        RECT 764.700 3.500 772.500 4.300 ;
        RECT 773.660 3.500 781.460 4.300 ;
        RECT 782.620 3.500 790.420 4.300 ;
        RECT 791.580 3.500 799.380 4.300 ;
        RECT 800.540 3.500 808.340 4.300 ;
        RECT 809.500 3.500 817.300 4.300 ;
        RECT 818.460 3.500 826.260 4.300 ;
        RECT 827.420 3.500 835.220 4.300 ;
        RECT 836.380 3.500 844.180 4.300 ;
        RECT 845.340 3.500 853.140 4.300 ;
        RECT 854.300 3.500 862.100 4.300 ;
        RECT 863.260 3.500 871.060 4.300 ;
        RECT 872.220 3.500 880.020 4.300 ;
        RECT 881.180 3.500 888.980 4.300 ;
        RECT 890.140 3.500 897.940 4.300 ;
        RECT 899.100 3.500 906.900 4.300 ;
        RECT 908.060 3.500 915.860 4.300 ;
        RECT 917.020 3.500 924.820 4.300 ;
        RECT 925.980 3.500 933.780 4.300 ;
        RECT 934.940 3.500 942.740 4.300 ;
        RECT 943.900 3.500 951.700 4.300 ;
        RECT 952.860 3.500 994.420 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 656.060 996.000 682.220 ;
        RECT 4.000 654.900 995.700 656.060 ;
        RECT 4.000 649.340 996.000 654.900 ;
        RECT 4.300 648.220 996.000 649.340 ;
        RECT 4.300 648.180 995.700 648.220 ;
        RECT 4.000 647.060 995.700 648.180 ;
        RECT 4.000 642.620 996.000 647.060 ;
        RECT 4.300 641.460 996.000 642.620 ;
        RECT 4.000 640.380 996.000 641.460 ;
        RECT 4.000 639.220 995.700 640.380 ;
        RECT 4.000 635.900 996.000 639.220 ;
        RECT 4.300 634.740 996.000 635.900 ;
        RECT 4.000 632.540 996.000 634.740 ;
        RECT 4.000 631.380 995.700 632.540 ;
        RECT 4.000 629.180 996.000 631.380 ;
        RECT 4.300 628.020 996.000 629.180 ;
        RECT 4.000 624.700 996.000 628.020 ;
        RECT 4.000 623.540 995.700 624.700 ;
        RECT 4.000 622.460 996.000 623.540 ;
        RECT 4.300 621.300 996.000 622.460 ;
        RECT 4.000 616.860 996.000 621.300 ;
        RECT 4.000 615.740 995.700 616.860 ;
        RECT 4.300 615.700 995.700 615.740 ;
        RECT 4.300 614.580 996.000 615.700 ;
        RECT 4.000 609.020 996.000 614.580 ;
        RECT 4.300 607.860 995.700 609.020 ;
        RECT 4.000 602.300 996.000 607.860 ;
        RECT 4.300 601.180 996.000 602.300 ;
        RECT 4.300 601.140 995.700 601.180 ;
        RECT 4.000 600.020 995.700 601.140 ;
        RECT 4.000 595.580 996.000 600.020 ;
        RECT 4.300 594.420 996.000 595.580 ;
        RECT 4.000 593.340 996.000 594.420 ;
        RECT 4.000 592.180 995.700 593.340 ;
        RECT 4.000 588.860 996.000 592.180 ;
        RECT 4.300 587.700 996.000 588.860 ;
        RECT 4.000 585.500 996.000 587.700 ;
        RECT 4.000 584.340 995.700 585.500 ;
        RECT 4.000 582.140 996.000 584.340 ;
        RECT 4.300 580.980 996.000 582.140 ;
        RECT 4.000 577.660 996.000 580.980 ;
        RECT 4.000 576.500 995.700 577.660 ;
        RECT 4.000 575.420 996.000 576.500 ;
        RECT 4.300 574.260 996.000 575.420 ;
        RECT 4.000 569.820 996.000 574.260 ;
        RECT 4.000 568.700 995.700 569.820 ;
        RECT 4.300 568.660 995.700 568.700 ;
        RECT 4.300 567.540 996.000 568.660 ;
        RECT 4.000 561.980 996.000 567.540 ;
        RECT 4.300 560.820 995.700 561.980 ;
        RECT 4.000 555.260 996.000 560.820 ;
        RECT 4.300 554.140 996.000 555.260 ;
        RECT 4.300 554.100 995.700 554.140 ;
        RECT 4.000 552.980 995.700 554.100 ;
        RECT 4.000 548.540 996.000 552.980 ;
        RECT 4.300 547.380 996.000 548.540 ;
        RECT 4.000 546.300 996.000 547.380 ;
        RECT 4.000 545.140 995.700 546.300 ;
        RECT 4.000 541.820 996.000 545.140 ;
        RECT 4.300 540.660 996.000 541.820 ;
        RECT 4.000 538.460 996.000 540.660 ;
        RECT 4.000 537.300 995.700 538.460 ;
        RECT 4.000 535.100 996.000 537.300 ;
        RECT 4.300 533.940 996.000 535.100 ;
        RECT 4.000 530.620 996.000 533.940 ;
        RECT 4.000 529.460 995.700 530.620 ;
        RECT 4.000 528.380 996.000 529.460 ;
        RECT 4.300 527.220 996.000 528.380 ;
        RECT 4.000 522.780 996.000 527.220 ;
        RECT 4.000 521.660 995.700 522.780 ;
        RECT 4.300 521.620 995.700 521.660 ;
        RECT 4.300 520.500 996.000 521.620 ;
        RECT 4.000 514.940 996.000 520.500 ;
        RECT 4.300 513.780 995.700 514.940 ;
        RECT 4.000 508.220 996.000 513.780 ;
        RECT 4.300 507.100 996.000 508.220 ;
        RECT 4.300 507.060 995.700 507.100 ;
        RECT 4.000 505.940 995.700 507.060 ;
        RECT 4.000 501.500 996.000 505.940 ;
        RECT 4.300 500.340 996.000 501.500 ;
        RECT 4.000 499.260 996.000 500.340 ;
        RECT 4.000 498.100 995.700 499.260 ;
        RECT 4.000 494.780 996.000 498.100 ;
        RECT 4.300 493.620 996.000 494.780 ;
        RECT 4.000 491.420 996.000 493.620 ;
        RECT 4.000 490.260 995.700 491.420 ;
        RECT 4.000 488.060 996.000 490.260 ;
        RECT 4.300 486.900 996.000 488.060 ;
        RECT 4.000 483.580 996.000 486.900 ;
        RECT 4.000 482.420 995.700 483.580 ;
        RECT 4.000 481.340 996.000 482.420 ;
        RECT 4.300 480.180 996.000 481.340 ;
        RECT 4.000 475.740 996.000 480.180 ;
        RECT 4.000 474.620 995.700 475.740 ;
        RECT 4.300 474.580 995.700 474.620 ;
        RECT 4.300 473.460 996.000 474.580 ;
        RECT 4.000 467.900 996.000 473.460 ;
        RECT 4.300 466.740 995.700 467.900 ;
        RECT 4.000 461.180 996.000 466.740 ;
        RECT 4.300 460.060 996.000 461.180 ;
        RECT 4.300 460.020 995.700 460.060 ;
        RECT 4.000 458.900 995.700 460.020 ;
        RECT 4.000 454.460 996.000 458.900 ;
        RECT 4.300 453.300 996.000 454.460 ;
        RECT 4.000 452.220 996.000 453.300 ;
        RECT 4.000 451.060 995.700 452.220 ;
        RECT 4.000 447.740 996.000 451.060 ;
        RECT 4.300 446.580 996.000 447.740 ;
        RECT 4.000 444.380 996.000 446.580 ;
        RECT 4.000 443.220 995.700 444.380 ;
        RECT 4.000 441.020 996.000 443.220 ;
        RECT 4.300 439.860 996.000 441.020 ;
        RECT 4.000 436.540 996.000 439.860 ;
        RECT 4.000 435.380 995.700 436.540 ;
        RECT 4.000 434.300 996.000 435.380 ;
        RECT 4.300 433.140 996.000 434.300 ;
        RECT 4.000 428.700 996.000 433.140 ;
        RECT 4.000 427.580 995.700 428.700 ;
        RECT 4.300 427.540 995.700 427.580 ;
        RECT 4.300 426.420 996.000 427.540 ;
        RECT 4.000 420.860 996.000 426.420 ;
        RECT 4.300 419.700 995.700 420.860 ;
        RECT 4.000 414.140 996.000 419.700 ;
        RECT 4.300 413.020 996.000 414.140 ;
        RECT 4.300 412.980 995.700 413.020 ;
        RECT 4.000 411.860 995.700 412.980 ;
        RECT 4.000 407.420 996.000 411.860 ;
        RECT 4.300 406.260 996.000 407.420 ;
        RECT 4.000 405.180 996.000 406.260 ;
        RECT 4.000 404.020 995.700 405.180 ;
        RECT 4.000 400.700 996.000 404.020 ;
        RECT 4.300 399.540 996.000 400.700 ;
        RECT 4.000 397.340 996.000 399.540 ;
        RECT 4.000 396.180 995.700 397.340 ;
        RECT 4.000 393.980 996.000 396.180 ;
        RECT 4.300 392.820 996.000 393.980 ;
        RECT 4.000 389.500 996.000 392.820 ;
        RECT 4.000 388.340 995.700 389.500 ;
        RECT 4.000 387.260 996.000 388.340 ;
        RECT 4.300 386.100 996.000 387.260 ;
        RECT 4.000 381.660 996.000 386.100 ;
        RECT 4.000 380.540 995.700 381.660 ;
        RECT 4.300 380.500 995.700 380.540 ;
        RECT 4.300 379.380 996.000 380.500 ;
        RECT 4.000 373.820 996.000 379.380 ;
        RECT 4.300 372.660 995.700 373.820 ;
        RECT 4.000 367.100 996.000 372.660 ;
        RECT 4.300 365.980 996.000 367.100 ;
        RECT 4.300 365.940 995.700 365.980 ;
        RECT 4.000 364.820 995.700 365.940 ;
        RECT 4.000 360.380 996.000 364.820 ;
        RECT 4.300 359.220 996.000 360.380 ;
        RECT 4.000 358.140 996.000 359.220 ;
        RECT 4.000 356.980 995.700 358.140 ;
        RECT 4.000 353.660 996.000 356.980 ;
        RECT 4.300 352.500 996.000 353.660 ;
        RECT 4.000 350.300 996.000 352.500 ;
        RECT 4.000 349.140 995.700 350.300 ;
        RECT 4.000 346.940 996.000 349.140 ;
        RECT 4.300 345.780 996.000 346.940 ;
        RECT 4.000 342.460 996.000 345.780 ;
        RECT 4.000 341.300 995.700 342.460 ;
        RECT 4.000 340.220 996.000 341.300 ;
        RECT 4.300 339.060 996.000 340.220 ;
        RECT 4.000 334.620 996.000 339.060 ;
        RECT 4.000 333.500 995.700 334.620 ;
        RECT 4.300 333.460 995.700 333.500 ;
        RECT 4.300 332.340 996.000 333.460 ;
        RECT 4.000 326.780 996.000 332.340 ;
        RECT 4.300 325.620 995.700 326.780 ;
        RECT 4.000 320.060 996.000 325.620 ;
        RECT 4.300 318.940 996.000 320.060 ;
        RECT 4.300 318.900 995.700 318.940 ;
        RECT 4.000 317.780 995.700 318.900 ;
        RECT 4.000 313.340 996.000 317.780 ;
        RECT 4.300 312.180 996.000 313.340 ;
        RECT 4.000 311.100 996.000 312.180 ;
        RECT 4.000 309.940 995.700 311.100 ;
        RECT 4.000 306.620 996.000 309.940 ;
        RECT 4.300 305.460 996.000 306.620 ;
        RECT 4.000 303.260 996.000 305.460 ;
        RECT 4.000 302.100 995.700 303.260 ;
        RECT 4.000 299.900 996.000 302.100 ;
        RECT 4.300 298.740 996.000 299.900 ;
        RECT 4.000 295.420 996.000 298.740 ;
        RECT 4.000 294.260 995.700 295.420 ;
        RECT 4.000 293.180 996.000 294.260 ;
        RECT 4.300 292.020 996.000 293.180 ;
        RECT 4.000 287.580 996.000 292.020 ;
        RECT 4.000 286.460 995.700 287.580 ;
        RECT 4.300 286.420 995.700 286.460 ;
        RECT 4.300 285.300 996.000 286.420 ;
        RECT 4.000 279.740 996.000 285.300 ;
        RECT 4.300 278.580 995.700 279.740 ;
        RECT 4.000 273.020 996.000 278.580 ;
        RECT 4.300 271.900 996.000 273.020 ;
        RECT 4.300 271.860 995.700 271.900 ;
        RECT 4.000 270.740 995.700 271.860 ;
        RECT 4.000 266.300 996.000 270.740 ;
        RECT 4.300 265.140 996.000 266.300 ;
        RECT 4.000 264.060 996.000 265.140 ;
        RECT 4.000 262.900 995.700 264.060 ;
        RECT 4.000 259.580 996.000 262.900 ;
        RECT 4.300 258.420 996.000 259.580 ;
        RECT 4.000 256.220 996.000 258.420 ;
        RECT 4.000 255.060 995.700 256.220 ;
        RECT 4.000 252.860 996.000 255.060 ;
        RECT 4.300 251.700 996.000 252.860 ;
        RECT 4.000 248.380 996.000 251.700 ;
        RECT 4.000 247.220 995.700 248.380 ;
        RECT 4.000 246.140 996.000 247.220 ;
        RECT 4.300 244.980 996.000 246.140 ;
        RECT 4.000 240.540 996.000 244.980 ;
        RECT 4.000 239.420 995.700 240.540 ;
        RECT 4.300 239.380 995.700 239.420 ;
        RECT 4.300 238.260 996.000 239.380 ;
        RECT 4.000 232.700 996.000 238.260 ;
        RECT 4.300 231.540 995.700 232.700 ;
        RECT 4.000 225.980 996.000 231.540 ;
        RECT 4.300 224.860 996.000 225.980 ;
        RECT 4.300 224.820 995.700 224.860 ;
        RECT 4.000 223.700 995.700 224.820 ;
        RECT 4.000 219.260 996.000 223.700 ;
        RECT 4.300 218.100 996.000 219.260 ;
        RECT 4.000 217.020 996.000 218.100 ;
        RECT 4.000 215.860 995.700 217.020 ;
        RECT 4.000 212.540 996.000 215.860 ;
        RECT 4.300 211.380 996.000 212.540 ;
        RECT 4.000 209.180 996.000 211.380 ;
        RECT 4.000 208.020 995.700 209.180 ;
        RECT 4.000 205.820 996.000 208.020 ;
        RECT 4.300 204.660 996.000 205.820 ;
        RECT 4.000 201.340 996.000 204.660 ;
        RECT 4.000 200.180 995.700 201.340 ;
        RECT 4.000 199.100 996.000 200.180 ;
        RECT 4.300 197.940 996.000 199.100 ;
        RECT 4.000 193.500 996.000 197.940 ;
        RECT 4.000 192.380 995.700 193.500 ;
        RECT 4.300 192.340 995.700 192.380 ;
        RECT 4.300 191.220 996.000 192.340 ;
        RECT 4.000 185.660 996.000 191.220 ;
        RECT 4.300 184.500 995.700 185.660 ;
        RECT 4.000 178.940 996.000 184.500 ;
        RECT 4.300 177.820 996.000 178.940 ;
        RECT 4.300 177.780 995.700 177.820 ;
        RECT 4.000 176.660 995.700 177.780 ;
        RECT 4.000 172.220 996.000 176.660 ;
        RECT 4.300 171.060 996.000 172.220 ;
        RECT 4.000 169.980 996.000 171.060 ;
        RECT 4.000 168.820 995.700 169.980 ;
        RECT 4.000 165.500 996.000 168.820 ;
        RECT 4.300 164.340 996.000 165.500 ;
        RECT 4.000 162.140 996.000 164.340 ;
        RECT 4.000 160.980 995.700 162.140 ;
        RECT 4.000 158.780 996.000 160.980 ;
        RECT 4.300 157.620 996.000 158.780 ;
        RECT 4.000 154.300 996.000 157.620 ;
        RECT 4.000 153.140 995.700 154.300 ;
        RECT 4.000 152.060 996.000 153.140 ;
        RECT 4.300 150.900 996.000 152.060 ;
        RECT 4.000 146.460 996.000 150.900 ;
        RECT 4.000 145.340 995.700 146.460 ;
        RECT 4.300 145.300 995.700 145.340 ;
        RECT 4.300 144.180 996.000 145.300 ;
        RECT 4.000 138.620 996.000 144.180 ;
        RECT 4.300 137.460 995.700 138.620 ;
        RECT 4.000 131.900 996.000 137.460 ;
        RECT 4.300 130.780 996.000 131.900 ;
        RECT 4.300 130.740 995.700 130.780 ;
        RECT 4.000 129.620 995.700 130.740 ;
        RECT 4.000 125.180 996.000 129.620 ;
        RECT 4.300 124.020 996.000 125.180 ;
        RECT 4.000 122.940 996.000 124.020 ;
        RECT 4.000 121.780 995.700 122.940 ;
        RECT 4.000 118.460 996.000 121.780 ;
        RECT 4.300 117.300 996.000 118.460 ;
        RECT 4.000 115.100 996.000 117.300 ;
        RECT 4.000 113.940 995.700 115.100 ;
        RECT 4.000 111.740 996.000 113.940 ;
        RECT 4.300 110.580 996.000 111.740 ;
        RECT 4.000 107.260 996.000 110.580 ;
        RECT 4.000 106.100 995.700 107.260 ;
        RECT 4.000 105.020 996.000 106.100 ;
        RECT 4.300 103.860 996.000 105.020 ;
        RECT 4.000 99.420 996.000 103.860 ;
        RECT 4.000 98.300 995.700 99.420 ;
        RECT 4.300 98.260 995.700 98.300 ;
        RECT 4.300 97.140 996.000 98.260 ;
        RECT 4.000 91.580 996.000 97.140 ;
        RECT 4.300 90.420 995.700 91.580 ;
        RECT 4.000 84.860 996.000 90.420 ;
        RECT 4.300 83.740 996.000 84.860 ;
        RECT 4.300 83.700 995.700 83.740 ;
        RECT 4.000 82.580 995.700 83.700 ;
        RECT 4.000 78.140 996.000 82.580 ;
        RECT 4.300 76.980 996.000 78.140 ;
        RECT 4.000 75.900 996.000 76.980 ;
        RECT 4.000 74.740 995.700 75.900 ;
        RECT 4.000 71.420 996.000 74.740 ;
        RECT 4.300 70.260 996.000 71.420 ;
        RECT 4.000 68.060 996.000 70.260 ;
        RECT 4.000 66.900 995.700 68.060 ;
        RECT 4.000 64.700 996.000 66.900 ;
        RECT 4.300 63.540 996.000 64.700 ;
        RECT 4.000 60.220 996.000 63.540 ;
        RECT 4.000 59.060 995.700 60.220 ;
        RECT 4.000 57.980 996.000 59.060 ;
        RECT 4.300 56.820 996.000 57.980 ;
        RECT 4.000 52.380 996.000 56.820 ;
        RECT 4.000 51.260 995.700 52.380 ;
        RECT 4.300 51.220 995.700 51.260 ;
        RECT 4.300 50.100 996.000 51.220 ;
        RECT 4.000 44.540 996.000 50.100 ;
        RECT 4.000 43.380 995.700 44.540 ;
        RECT 4.000 12.460 996.000 43.380 ;
      LAYER Metal4 ;
        RECT 158.060 34.250 175.540 671.350 ;
        RECT 177.740 34.250 252.340 671.350 ;
        RECT 254.540 34.250 329.140 671.350 ;
        RECT 331.340 34.250 405.940 671.350 ;
        RECT 408.140 34.250 482.740 671.350 ;
        RECT 484.940 34.250 559.540 671.350 ;
        RECT 561.740 34.250 636.340 671.350 ;
        RECT 638.540 34.250 713.140 671.350 ;
        RECT 715.340 34.250 789.940 671.350 ;
        RECT 792.140 34.250 866.740 671.350 ;
        RECT 868.940 34.250 943.540 671.350 ;
        RECT 945.740 34.250 954.660 671.350 ;
  END
END wrapped_as2650
END LIBRARY

