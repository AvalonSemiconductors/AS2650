VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO timers
  CLASS BLOCK ;
  FOREIGN timers ;
  ORIGIN 0.000 0.000 ;
  SIZE 425.000 BY 425.000 ;
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.680 4.000 16.240 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.920 4.000 46.480 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 76.160 4.000 76.720 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.400 4.000 106.960 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 136.640 4.000 137.200 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.880 4.000 167.440 ;
    END
  END addr[5]
  PIN bus_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END bus_cyc
  PIN bus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END bus_we
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 197.120 4.000 197.680 ;
    END
  END data_in[0]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 227.360 4.000 227.920 ;
    END
  END data_in[1]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.600 4.000 258.160 ;
    END
  END data_in[2]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 287.840 4.000 288.400 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.080 4.000 318.640 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 348.320 4.000 348.880 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 378.560 4.000 379.120 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 408.800 4.000 409.360 ;
    END
  END data_in[7]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 421.000 28.000 425.000 28.560 ;
    END
  END data_out[0]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 421.000 80.640 425.000 81.200 ;
    END
  END data_out[1]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 421.000 133.280 425.000 133.840 ;
    END
  END data_out[2]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 421.000 185.920 425.000 186.480 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 421.000 238.560 425.000 239.120 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 421.000 291.200 425.000 291.760 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 421.000 343.840 425.000 344.400 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 421.000 396.480 425.000 397.040 ;
    END
  END data_out[7]
  PIN irq1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 4.000 ;
    END
  END irq1
  PIN irq2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END irq2
  PIN irq5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END irq5
  PIN pwm0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 421.000 212.240 425.000 ;
    END
  END pwm0
  PIN pwm1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 421.000 297.360 425.000 ;
    END
  END pwm1
  PIN pwm2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 381.920 421.000 382.480 425.000 ;
    END
  END pwm2
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 0.000 306.320 4.000 ;
    END
  END rst
  PIN tmr0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 0.000 353.360 4.000 ;
    END
  END tmr0_clk
  PIN tmr0_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 421.000 42.000 425.000 ;
    END
  END tmr0_o
  PIN tmr1_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 0.000 400.400 4.000 ;
    END
  END tmr1_clk
  PIN tmr1_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 421.000 127.120 425.000 ;
    END
  END tmr1_o
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 407.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 407.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 407.980 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 407.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 407.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 407.980 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 0.000 259.280 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 417.760 407.980 ;
      LAYER Metal2 ;
        RECT 5.740 420.700 41.140 421.000 ;
        RECT 42.300 420.700 126.260 421.000 ;
        RECT 127.420 420.700 211.380 421.000 ;
        RECT 212.540 420.700 296.500 421.000 ;
        RECT 297.660 420.700 381.620 421.000 ;
        RECT 382.780 420.700 415.940 421.000 ;
        RECT 5.740 4.300 415.940 420.700 ;
        RECT 5.740 4.000 23.220 4.300 ;
        RECT 24.380 4.000 70.260 4.300 ;
        RECT 71.420 4.000 117.300 4.300 ;
        RECT 118.460 4.000 164.340 4.300 ;
        RECT 165.500 4.000 211.380 4.300 ;
        RECT 212.540 4.000 258.420 4.300 ;
        RECT 259.580 4.000 305.460 4.300 ;
        RECT 306.620 4.000 352.500 4.300 ;
        RECT 353.660 4.000 399.540 4.300 ;
        RECT 400.700 4.000 415.940 4.300 ;
      LAYER Metal3 ;
        RECT 4.300 408.500 421.000 409.220 ;
        RECT 4.000 397.340 421.000 408.500 ;
        RECT 4.000 396.180 420.700 397.340 ;
        RECT 4.000 379.420 421.000 396.180 ;
        RECT 4.300 378.260 421.000 379.420 ;
        RECT 4.000 349.180 421.000 378.260 ;
        RECT 4.300 348.020 421.000 349.180 ;
        RECT 4.000 344.700 421.000 348.020 ;
        RECT 4.000 343.540 420.700 344.700 ;
        RECT 4.000 318.940 421.000 343.540 ;
        RECT 4.300 317.780 421.000 318.940 ;
        RECT 4.000 292.060 421.000 317.780 ;
        RECT 4.000 290.900 420.700 292.060 ;
        RECT 4.000 288.700 421.000 290.900 ;
        RECT 4.300 287.540 421.000 288.700 ;
        RECT 4.000 258.460 421.000 287.540 ;
        RECT 4.300 257.300 421.000 258.460 ;
        RECT 4.000 239.420 421.000 257.300 ;
        RECT 4.000 238.260 420.700 239.420 ;
        RECT 4.000 228.220 421.000 238.260 ;
        RECT 4.300 227.060 421.000 228.220 ;
        RECT 4.000 197.980 421.000 227.060 ;
        RECT 4.300 196.820 421.000 197.980 ;
        RECT 4.000 186.780 421.000 196.820 ;
        RECT 4.000 185.620 420.700 186.780 ;
        RECT 4.000 167.740 421.000 185.620 ;
        RECT 4.300 166.580 421.000 167.740 ;
        RECT 4.000 137.500 421.000 166.580 ;
        RECT 4.300 136.340 421.000 137.500 ;
        RECT 4.000 134.140 421.000 136.340 ;
        RECT 4.000 132.980 420.700 134.140 ;
        RECT 4.000 107.260 421.000 132.980 ;
        RECT 4.300 106.100 421.000 107.260 ;
        RECT 4.000 81.500 421.000 106.100 ;
        RECT 4.000 80.340 420.700 81.500 ;
        RECT 4.000 77.020 421.000 80.340 ;
        RECT 4.300 75.860 421.000 77.020 ;
        RECT 4.000 46.780 421.000 75.860 ;
        RECT 4.300 45.620 421.000 46.780 ;
        RECT 4.000 28.860 421.000 45.620 ;
        RECT 4.000 27.700 420.700 28.860 ;
        RECT 4.000 16.540 421.000 27.700 ;
        RECT 4.300 15.540 421.000 16.540 ;
      LAYER Metal4 ;
        RECT 26.460 25.850 98.740 370.630 ;
        RECT 100.940 25.850 175.540 370.630 ;
        RECT 177.740 25.850 252.340 370.630 ;
        RECT 254.540 25.850 329.140 370.630 ;
        RECT 331.340 25.850 390.180 370.630 ;
  END
END timers
END LIBRARY

