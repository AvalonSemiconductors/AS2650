// This is the unpowered netlist.
module gpios (RXD,
    TXD,
    bus_cyc,
    bus_we,
    irq0,
    irq6,
    irq7,
    pwm0,
    pwm1,
    pwm2,
    rst,
    tmr0_clk,
    tmr0_o,
    tmr1_clk,
    tmr1_o,
    wb_clk_i,
    addr,
    data_in,
    data_out,
    io_in,
    io_oeb,
    io_out,
    la_data_out);
 output RXD;
 input TXD;
 input bus_cyc;
 input bus_we;
 output irq0;
 output irq6;
 output irq7;
 input pwm0;
 input pwm1;
 input pwm2;
 input rst;
 output tmr0_clk;
 input tmr0_o;
 output tmr1_clk;
 input tmr1_o;
 input wb_clk_i;
 input [3:0] addr;
 input [7:0] data_in;
 output [7:0] data_out;
 input [15:0] io_in;
 output [15:0] io_oeb;
 output [15:0] io_out;
 output [7:0] la_data_out;

 wire \DDRA[0] ;
 wire \DDRA[1] ;
 wire \DDRA[2] ;
 wire \DDRA[3] ;
 wire \DDRA[4] ;
 wire \DDRA[5] ;
 wire \DDRA[6] ;
 wire \DDRA[7] ;
 wire \DDRB[0] ;
 wire \DDRB[1] ;
 wire \DDRB[2] ;
 wire \DDRB[3] ;
 wire \DDRB[4] ;
 wire \DDRB[5] ;
 wire \DDRB[6] ;
 wire \DDRB[7] ;
 wire \PORTA[0] ;
 wire \PORTA[1] ;
 wire \PORTA[2] ;
 wire \PORTA[3] ;
 wire \PORTA[4] ;
 wire \PORTA[5] ;
 wire \PORTA[6] ;
 wire \PORTA[7] ;
 wire \PORTB[0] ;
 wire \PORTB[1] ;
 wire \PORTB[2] ;
 wire \PORTB[3] ;
 wire \PORTB[4] ;
 wire \PORTB[5] ;
 wire \PORTB[6] ;
 wire \PORTB[7] ;
 wire \SPA[0] ;
 wire \SPA[1] ;
 wire \SPA[2] ;
 wire \SPA[3] ;
 wire \SPA[4] ;
 wire \SPA[5] ;
 wire \SPA[6] ;
 wire \SPA[7] ;
 wire \SPB[0] ;
 wire \SPB[1] ;
 wire \SPB[2] ;
 wire \SPB[3] ;
 wire \SPB[4] ;
 wire \SPB[5] ;
 wire \SPB[6] ;
 wire \SPB[7] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire last_irg6_trigger;
 wire last_irq0_trigger;
 wire last_irq7_trigger;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__398__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__400__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__400__S (.I(\SPA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__I1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__S (.I(\SPA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__I0 (.I(\PORTA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__I1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__S (.I(\SPA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__409__I1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__409__S (.I(\SPA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__411__I0 (.I(\PORTA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__411__S (.I(\SPA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__I (.I(\SPA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__A1 (.I(_079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__416__A1 (.I(\SPA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__417__A1 (.I(\SPA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__418__A1 (.I(\SPA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__418__A2 (.I(\DDRA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__A1 (.I(\SPA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__A1 (.I(\SPA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__425__I (.I(_083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__426__I0 (.I(\PORTB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__426__S (.I(\SPB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__428__I (.I(\SPB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__430__I (.I(_086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__431__I (.I(\SPB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__432__A1 (.I(_087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__435__A2 (.I(\PORTB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__A1 (.I(_091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__A2 (.I(\PORTB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__440__I (.I(\SPB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__A1 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__A2 (.I(\PORTB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__443__I (.I(\SPB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__444__A1 (.I(_095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__A1 (.I(\SPB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__A2 (.I(\DDRA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__A2 (.I(\DDRA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__449__A1 (.I(_079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__450__A2 (.I(\DDRB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__A2 (.I(\DDRB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__452__A1 (.I(_087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__452__A2 (.I(\DDRB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__453__A2 (.I(\DDRB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__454__A1 (.I(_091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__454__A2 (.I(\DDRB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__A1 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__A2 (.I(\DDRB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__456__A1 (.I(_095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__456__A2 (.I(\DDRB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__A1 (.I(\SPB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__A2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__459__A1 (.I(\SPB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__461__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__I (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__A1 (.I(\SPA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__A2 (.I(_102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__475__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__B2 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__C2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__493__I (.I(_129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__494__A1 (.I(\DDRB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__500__I (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__I (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__I (.I(_141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__B2 (.I(\DDRA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__C (.I(_148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__A1 (.I(_150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__518__I (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__I (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__A2 (.I(_141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__C1 (.I(\SPA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__I (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__A1 (.I(\SPB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__B2 (.I(\PORTB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__C (.I(_148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__528__A1 (.I(\SPB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__A1 (.I(\DDRB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__B2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__532__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__B2 (.I(\DDRA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__A1 (.I(\SPB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__B2 (.I(\DDRB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__541__A2 (.I(_141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__541__C1 (.I(\SPA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__542__I (.I(_129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__545__A1 (.I(_150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__A1 (.I(\DDRB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__549__A1 (.I(\PORTB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__549__B2 (.I(\DDRA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__551__B2 (.I(\PORTA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__551__C1 (.I(\SPA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__556__B2 (.I(\DDRB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__A2 (.I(_141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__B1 (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__C1 (.I(\SPA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__558__A1 (.I(\PORTB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__560__A1 (.I(_150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__563__A1 (.I(\DDRB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__563__C2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__B2 (.I(\PORTA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__C1 (.I(\SPA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__565__A1 (.I(\SPB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__566__A1 (.I(\PORTB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__566__B2 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__568__C (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__572__A1 (.I(_200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__572__B (.I(_150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__572__C (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__573__A1 (.I(\DDRB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__573__B2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__574__B2 (.I(\SPA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__575__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__576__A1 (.I(\SPB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__578__C (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__583__A1 (.I(_208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__583__A3 (.I(_211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__584__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__A2 (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__586__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__589__A3 (.I(_211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__590__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__591__A2 (.I(_218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__592__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__596__A1 (.I(_222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__596__A3 (.I(_211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__597__A2 (.I(_102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__598__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__599__A1 (.I(_221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__602__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__602__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__604__I (.I(_229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__605__A1 (.I(_226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__607__A2 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__611__I (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__614__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__615__C (.I(_221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__616__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__617__A1 (.I(_240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__622__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__623__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__625__C (.I(_247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__626__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__627__A1 (.I(_248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__631__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__632__C (.I(_247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__633__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__634__A1 (.I(_253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__638__A1 (.I(_256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__638__A2 (.I(_229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__640__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__642__B (.I(_260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__644__A2 (.I(_261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__646__A1 (.I(_226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__647__A2 (.I(_211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__649__A1 (.I(\DDRA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__650__B (.I(_260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__651__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__652__A1 (.I(_268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__654__B (.I(_260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__655__A1 (.I(_240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__656__A1 (.I(\DDRA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__657__B (.I(_260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__658__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__659__A1 (.I(_273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__664__A1 (.I(_248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__666__A1 (.I(\DDRA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__668__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__669__A1 (.I(_281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__672__A1 (.I(_253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__675__A1 (.I(_256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__681__I (.I(_290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__682__A1 (.I(_226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__685__A1 (.I(\DDRB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__688__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__689__C (.I(_247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__690__A1 (.I(_240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__691__A1 (.I(\DDRB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__693__A1 (.I(_273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__694__A1 (.I(\DDRB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__696__A1 (.I(_248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__698__A1 (.I(\DDRB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__701__A1 (.I(_281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__701__A2 (.I(_290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__702__A1 (.I(\DDRB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__704__A1 (.I(_253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__704__A2 (.I(_290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__705__A1 (.I(\DDRB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__707__A1 (.I(_256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__707__A2 (.I(_290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__708__A1 (.I(\DDRB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__710__A1 (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__710__A2 (.I(_261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__712__A1 (.I(_226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__713__A2 (.I(_261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__716__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__719__A1 (.I(_268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__722__A1 (.I(_240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__725__A1 (.I(_273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__729__A1 (.I(_248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__731__A1 (.I(\PORTA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__734__A1 (.I(_281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__737__A1 (.I(_253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__738__A1 (.I(\PORTA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__740__A1 (.I(_256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__743__A1 (.I(_129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__743__A2 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__745__A1 (.I(_208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__746__A1 (.I(_129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__746__A2 (.I(_261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__751__A1 (.I(_268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__752__A1 (.I(\PORTB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__754__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__757__A1 (.I(_273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__761__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__763__A1 (.I(\PORTB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__766__A1 (.I(_281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__767__A1 (.I(\PORTB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__770__A1 (.I(\PORTB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__772__A1 (.I(_222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__775__A1 (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__778__A1 (.I(_208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__779__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__779__C (.I(_247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__780__A1 (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__780__A2 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__782__A1 (.I(_268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__783__A1 (.I(\SPA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__786__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__788__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__789__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__791__A1 (.I(\SPA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__793__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__794__A1 (.I(\SPA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__796__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__797__A1 (.I(\SPA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__800__A1 (.I(\SPA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__802__A1 (.I(_222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__803__A1 (.I(_079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__804__A1 (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__804__A2 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__807__A1 (.I(_208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__809__I (.I(\SPB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__810__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__812__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__815__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__816__A1 (.I(_087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__819__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__821__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__822__A1 (.I(_091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__824__A1 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__824__C (.I(_148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__825__A1 (.I(_222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__826__A1 (.I(_095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__826__C (.I(_148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__827__A1 (.I(_221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__827__A2 (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__828__A1 (.I(_221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__828__A2 (.I(_218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__829__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__831__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__838__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__839__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__840__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__841__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__843__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__844__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__845__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__846__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__847__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__848__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__849__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__850__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__851__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__852__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__853__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__854__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__855__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__865__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__866__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__867__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__868__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__873__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__875__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__877__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__879__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__880__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__888__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__889__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__890__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__891__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__892__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__893__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__894__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__895__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__896__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__897__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__898__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(data_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(data_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(data_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(data_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(data_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(data_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(TXD));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(pwm0));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(pwm1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(pwm2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(tmr0_o));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(tmr1_o));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(bus_cyc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(bus_we));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(data_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(data_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output48_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output79_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output80_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output81_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_152 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _397_ (.I(\SPA[0] ),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _398_ (.A1(_070_),
    .A2(\PORTA[0] ),
    .Z(_071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _399_ (.I(_071_),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _400_ (.I0(\PORTA[1] ),
    .I1(net1),
    .S(\SPA[1] ),
    .Z(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _401_ (.I(_072_),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _402_ (.I(\SPA[2] ),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _403_ (.A1(_073_),
    .A2(\PORTA[2] ),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _404_ (.I(_074_),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _405_ (.I0(\PORTA[3] ),
    .I1(net36),
    .S(\SPA[3] ),
    .Z(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _406_ (.I(_075_),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _407_ (.I0(\PORTA[4] ),
    .I1(net37),
    .S(\SPA[4] ),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _408_ (.I(_076_),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _409_ (.I0(\PORTA[5] ),
    .I1(net32),
    .S(\SPA[5] ),
    .Z(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _410_ (.I(_077_),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _411_ (.I0(\PORTA[6] ),
    .I1(net33),
    .S(\SPA[6] ),
    .Z(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _412_ (.I(_078_),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _413_ (.I(\SPA[7] ),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _414_ (.A1(_079_),
    .A2(\PORTA[7] ),
    .Z(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _415_ (.I(_080_),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _416_ (.A1(\SPA[1] ),
    .A2(\DDRA[1] ),
    .ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _417_ (.A1(\SPA[3] ),
    .A2(\DDRA[3] ),
    .ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _418_ (.A1(\SPA[4] ),
    .A2(\DDRA[4] ),
    .ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _419_ (.A1(\SPA[5] ),
    .A2(\DDRA[5] ),
    .ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _420_ (.A1(\SPA[6] ),
    .A2(\DDRA[6] ),
    .ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _421_ (.A1(_073_),
    .A2(net24),
    .Z(_081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _422_ (.I(_081_),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _423_ (.I(\SPB[0] ),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _424_ (.A1(_082_),
    .A2(\PORTB[0] ),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _425_ (.I(_083_),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _426_ (.I0(\PORTB[1] ),
    .I1(net34),
    .S(\SPB[1] ),
    .Z(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _427_ (.I(_084_),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _428_ (.I(\SPB[2] ),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _429_ (.A1(_085_),
    .A2(\PORTB[2] ),
    .Z(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _430_ (.I(_086_),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _431_ (.I(\SPB[3] ),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _432_ (.A1(_087_),
    .A2(\PORTB[3] ),
    .Z(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _433_ (.I(_088_),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _434_ (.I(\SPB[4] ),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _435_ (.A1(_089_),
    .A2(\PORTB[4] ),
    .Z(_090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _436_ (.I(_090_),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _437_ (.I(\SPB[5] ),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _438_ (.A1(_091_),
    .A2(\PORTB[5] ),
    .Z(_092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _439_ (.I(_092_),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _440_ (.I(\SPB[6] ),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _441_ (.A1(_093_),
    .A2(\PORTB[6] ),
    .Z(_094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _442_ (.I(_094_),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _443_ (.I(\SPB[7] ),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _444_ (.A1(_095_),
    .A2(\PORTB[7] ),
    .Z(_096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _445_ (.I(_096_),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _446_ (.A1(\SPB[1] ),
    .A2(\DDRB[1] ),
    .ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _447_ (.A1(_070_),
    .A2(\DDRA[0] ),
    .ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _448_ (.A1(_073_),
    .A2(\DDRA[2] ),
    .ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _449_ (.A1(_079_),
    .A2(\DDRA[7] ),
    .ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _450_ (.A1(_082_),
    .A2(\DDRB[0] ),
    .ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _451_ (.A1(_085_),
    .A2(\DDRB[2] ),
    .ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _452_ (.A1(_087_),
    .A2(\DDRB[3] ),
    .ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _453_ (.A1(_089_),
    .A2(\DDRB[4] ),
    .ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _454_ (.A1(_091_),
    .A2(\DDRB[5] ),
    .ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _455_ (.A1(_093_),
    .A2(\DDRB[6] ),
    .ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _456_ (.A1(_095_),
    .A2(\DDRB[7] ),
    .ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _457_ (.A1(\SPB[2] ),
    .A2(net17),
    .Z(_097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _458_ (.I(_097_),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _459_ (.A1(\SPB[3] ),
    .A2(net18),
    .Z(_098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _460_ (.I(_098_),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _461_ (.I(net35),
    .Z(_099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _462_ (.I(_099_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _463_ (.I(_100_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _464_ (.A1(\SPA[7] ),
    .A2(net29),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _465_ (.A1(_101_),
    .A2(_102_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _466_ (.I(net6),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _467_ (.I(_103_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _468_ (.I(_104_),
    .Z(_105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _469_ (.I(net39),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _470_ (.I(net5),
    .Z(_107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _471_ (.I(net3),
    .Z(_108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _472_ (.I(net4),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _473_ (.A1(net2),
    .A2(_108_),
    .A3(_109_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _474_ (.A1(_107_),
    .A2(_110_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _475_ (.I(_111_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _476_ (.I(net2),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _477_ (.I(_113_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _478_ (.I(net3),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _479_ (.I(_115_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _480_ (.I(net4),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _481_ (.I(_117_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _482_ (.I(net5),
    .Z(_119_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _483_ (.A1(_114_),
    .A2(_116_),
    .A3(_118_),
    .A4(_119_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _484_ (.I(_120_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _485_ (.I(_108_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _486_ (.A1(_114_),
    .A2(_122_),
    .A3(_118_),
    .A4(_119_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _487_ (.I(_123_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _488_ (.A1(\SPB[0] ),
    .A2(_112_),
    .B1(_121_),
    .B2(net79),
    .C1(_124_),
    .C2(net16),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _489_ (.A1(net4),
    .A2(net5),
    .Z(_126_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _490_ (.A1(_114_),
    .A2(_122_),
    .A3(_126_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _491_ (.I(_127_),
    .Z(_128_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _492_ (.A1(_113_),
    .A2(_116_),
    .A3(_126_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _493_ (.I(_129_),
    .Z(_130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _494_ (.A1(\DDRB[0] ),
    .A2(_128_),
    .B1(_130_),
    .B2(\PORTB[0] ),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _495_ (.I(_107_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _496_ (.A1(_113_),
    .A2(_108_),
    .A3(_109_),
    .A4(_132_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _497_ (.I(_133_),
    .Z(_134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _498_ (.I(net2),
    .Z(_135_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _499_ (.A1(_135_),
    .A2(_115_),
    .A3(_126_),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _500_ (.I(_136_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _501_ (.A1(net2),
    .A2(_108_),
    .A3(_117_),
    .A4(_107_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _502_ (.I(_138_),
    .Z(_139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _503_ (.A1(net82),
    .A2(_134_),
    .B1(_137_),
    .B2(\PORTA[0] ),
    .C1(\SPA[0] ),
    .C2(_139_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _504_ (.A1(_135_),
    .A2(_115_),
    .A3(_117_),
    .A4(_107_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _505_ (.I(_141_),
    .Z(_142_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _506_ (.A1(_132_),
    .A2(_110_),
    .Z(_143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _507_ (.I(_143_),
    .Z(_144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _508_ (.I(_103_),
    .Z(_145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _509_ (.A1(net30),
    .A2(_142_),
    .B1(_144_),
    .B2(\DDRA[0] ),
    .C(_145_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _510_ (.A1(_131_),
    .A2(_140_),
    .A3(_146_),
    .Z(_147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _511_ (.I(_099_),
    .Z(_148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _512_ (.A1(_105_),
    .A2(_106_),
    .B1(_125_),
    .B2(_147_),
    .C(_148_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _513_ (.I(net40),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _514_ (.A1(_122_),
    .A2(_109_),
    .B(_119_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _515_ (.I(_143_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _516_ (.A1(\DDRB[1] ),
    .A2(_128_),
    .B1(_151_),
    .B2(\DDRA[1] ),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _517_ (.A1(_150_),
    .A2(_152_),
    .Z(_153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _518_ (.I(_136_),
    .Z(_154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _519_ (.I(_138_),
    .Z(_155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _520_ (.A1(net31),
    .A2(_141_),
    .B1(_154_),
    .B2(\PORTA[1] ),
    .C1(\SPA[1] ),
    .C2(_155_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _521_ (.I(_123_),
    .Z(_157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _522_ (.A1(net83),
    .A2(_134_),
    .B1(_157_),
    .B2(net23),
    .C(_145_),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _523_ (.I(_111_),
    .Z(_159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _524_ (.A1(\SPB[1] ),
    .A2(_159_),
    .B1(_130_),
    .B2(\PORTB[1] ),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _525_ (.A1(_156_),
    .A2(_158_),
    .A3(_160_),
    .Z(_161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _526_ (.A1(_105_),
    .A2(_149_),
    .B1(_153_),
    .B2(_161_),
    .C(_148_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _527_ (.I(net41),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _528_ (.A1(\SPB[2] ),
    .A2(_112_),
    .B1(_130_),
    .B2(\PORTB[2] ),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _529_ (.A1(\DDRB[2] ),
    .A2(_128_),
    .B1(_124_),
    .B2(net24),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _530_ (.A1(_163_),
    .A2(_164_),
    .Z(_165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _531_ (.I(_133_),
    .Z(_166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _532_ (.A1(net17),
    .A2(_142_),
    .B1(_166_),
    .B2(net84),
    .C1(\SPA[2] ),
    .C2(_139_),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _533_ (.A1(\PORTA[2] ),
    .A2(_137_),
    .B1(_144_),
    .B2(\DDRA[2] ),
    .C(_145_),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _534_ (.A1(_167_),
    .A2(_168_),
    .Z(_169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _535_ (.I(_099_),
    .Z(_170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _536_ (.A1(_105_),
    .A2(_162_),
    .B1(_165_),
    .B2(_169_),
    .C(_170_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _537_ (.I(_104_),
    .Z(_171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _538_ (.I(net42),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _539_ (.I(_127_),
    .Z(_173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _540_ (.A1(\SPB[3] ),
    .A2(_112_),
    .B1(_173_),
    .B2(\DDRB[3] ),
    .C1(_151_),
    .C2(\DDRA[3] ),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _541_ (.A1(net18),
    .A2(_141_),
    .B1(_154_),
    .B2(\PORTA[3] ),
    .C1(\SPA[3] ),
    .C2(_155_),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _542_ (.I(_129_),
    .Z(_176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _543_ (.A1(\PORTB[3] ),
    .A2(_176_),
    .B1(_157_),
    .B2(net25),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _544_ (.A1(net85),
    .A2(_166_),
    .B(_104_),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _545_ (.A1(_150_),
    .A2(_175_),
    .A3(_177_),
    .A4(_178_),
    .Z(_179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _546_ (.A1(_171_),
    .A2(_172_),
    .B1(_174_),
    .B2(_179_),
    .C(_170_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _547_ (.I(net43),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _548_ (.A1(\DDRB[4] ),
    .A2(_128_),
    .B1(_157_),
    .B2(net26),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _549_ (.A1(\PORTB[4] ),
    .A2(_130_),
    .B1(_144_),
    .B2(\DDRA[4] ),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _550_ (.A1(_181_),
    .A2(_182_),
    .Z(_183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _551_ (.A1(net86),
    .A2(_134_),
    .B1(_137_),
    .B2(\PORTA[4] ),
    .C1(\SPA[4] ),
    .C2(_139_),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _552_ (.A1(\SPB[4] ),
    .A2(_159_),
    .B1(_142_),
    .B2(net19),
    .C(_145_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _553_ (.A1(_184_),
    .A2(_185_),
    .Z(_186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _554_ (.A1(_171_),
    .A2(_180_),
    .B1(_183_),
    .B2(_186_),
    .C(_170_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _555_ (.I(net44),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _556_ (.A1(\SPB[5] ),
    .A2(_112_),
    .B1(_173_),
    .B2(\DDRB[5] ),
    .C1(_151_),
    .C2(\DDRA[5] ),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _557_ (.A1(net20),
    .A2(_141_),
    .B1(_136_),
    .B2(\PORTA[5] ),
    .C1(\SPA[5] ),
    .C2(_155_),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _558_ (.A1(\PORTB[5] ),
    .A2(_176_),
    .B1(_157_),
    .B2(net27),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _559_ (.A1(net87),
    .A2(_166_),
    .B(_104_),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _560_ (.A1(_150_),
    .A2(_189_),
    .A3(_190_),
    .A4(_191_),
    .Z(_192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _561_ (.A1(_171_),
    .A2(_187_),
    .B1(_188_),
    .B2(_192_),
    .C(_170_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _562_ (.I(net45),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _563_ (.A1(\DDRB[6] ),
    .A2(_173_),
    .B1(_151_),
    .B2(\DDRA[6] ),
    .C1(_124_),
    .C2(net28),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _564_ (.A1(net88),
    .A2(_134_),
    .B1(_154_),
    .B2(\PORTA[6] ),
    .C1(\SPA[6] ),
    .C2(_155_),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _565_ (.A1(\SPB[6] ),
    .A2(_159_),
    .B1(_142_),
    .B2(net21),
    .C(_103_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _566_ (.A1(\PORTB[6] ),
    .A2(_176_),
    .B1(_120_),
    .B2(net80),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _567_ (.A1(_195_),
    .A2(_196_),
    .A3(_197_),
    .Z(_198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _568_ (.A1(_171_),
    .A2(_193_),
    .B1(_194_),
    .B2(_198_),
    .C(_100_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _569_ (.I(net46),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _570_ (.I(net22),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _571_ (.A1(_114_),
    .A2(_122_),
    .A3(_109_),
    .A4(_132_),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _572_ (.A1(_200_),
    .A2(_201_),
    .B(_150_),
    .C(net6),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _573_ (.A1(\DDRB[7] ),
    .A2(_173_),
    .B1(_124_),
    .B2(net29),
    .C(_202_),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _574_ (.A1(net89),
    .A2(_166_),
    .B1(_139_),
    .B2(\SPA[7] ),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _575_ (.A1(net81),
    .A2(_120_),
    .B1(_144_),
    .B2(\DDRA[7] ),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _576_ (.A1(\SPB[7] ),
    .A2(_159_),
    .B1(_176_),
    .B2(\PORTB[7] ),
    .C1(_137_),
    .C2(\PORTA[7] ),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _577_ (.A1(_204_),
    .A2(_205_),
    .A3(_206_),
    .Z(_207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _578_ (.A1(_199_),
    .A2(_105_),
    .B1(_203_),
    .B2(_207_),
    .C(_100_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _579_ (.I(net8),
    .Z(_208_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _580_ (.A1(net6),
    .A2(net7),
    .Z(_209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _581_ (.I(_209_),
    .Z(_210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _582_ (.I(_210_),
    .Z(_211_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _583_ (.A1(_208_),
    .A2(_121_),
    .A3(_211_),
    .ZN(_212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _584_ (.A1(\SPA[0] ),
    .A2(net16),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _585_ (.A1(last_irq0_trigger),
    .A2(_213_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _586_ (.A1(net79),
    .A2(_212_),
    .B(_214_),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _587_ (.A1(_101_),
    .A2(_215_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _588_ (.I(net14),
    .Z(_216_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _589_ (.A1(_216_),
    .A2(_121_),
    .A3(_211_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _590_ (.A1(\SPB[0] ),
    .A2(net30),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _591_ (.A1(last_irg6_trigger),
    .A2(_218_),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _592_ (.A1(net80),
    .A2(_217_),
    .B(_219_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _593_ (.A1(_101_),
    .A2(_220_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _594_ (.I(_099_),
    .Z(_221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _595_ (.I(net15),
    .Z(_222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _596_ (.A1(_222_),
    .A2(_121_),
    .A3(_211_),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _597_ (.A1(last_irq7_trigger),
    .A2(_102_),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _598_ (.A1(net81),
    .A2(_223_),
    .B(_224_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _599_ (.A1(_221_),
    .A2(_225_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _600_ (.I(net8),
    .Z(_226_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _601_ (.A1(_135_),
    .A2(_116_),
    .A3(_118_),
    .A4(_119_),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _602_ (.A1(net6),
    .A2(net7),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _603_ (.A1(_227_),
    .A2(_228_),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _604_ (.I(_229_),
    .Z(_230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _605_ (.A1(_226_),
    .A2(_230_),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _606_ (.I(_209_),
    .Z(_232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _607_ (.A1(_133_),
    .A2(_232_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _608_ (.I(_233_),
    .Z(_234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _609_ (.I(_234_),
    .Z(_235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _610_ (.A1(net82),
    .A2(_235_),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _611_ (.I(_100_),
    .Z(_237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _612_ (.A1(_231_),
    .A2(_236_),
    .B(_237_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _613_ (.I(net83),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _614_ (.A1(net9),
    .A2(_234_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _615_ (.A1(_238_),
    .A2(_235_),
    .B(_239_),
    .C(_221_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _616_ (.I(net10),
    .Z(_240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _617_ (.A1(_240_),
    .A2(_230_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _618_ (.I(_233_),
    .Z(_242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _619_ (.A1(net84),
    .A2(_242_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _620_ (.A1(_241_),
    .A2(_243_),
    .B(_237_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _621_ (.I(net85),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _622_ (.A1(net11),
    .A2(_234_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _623_ (.I(net35),
    .Z(_246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _624_ (.I(_246_),
    .Z(_247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _625_ (.A1(_244_),
    .A2(_235_),
    .B(_245_),
    .C(_247_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _626_ (.I(net12),
    .Z(_248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _627_ (.A1(_248_),
    .A2(_230_),
    .ZN(_249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _628_ (.A1(net86),
    .A2(_242_),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _629_ (.A1(_249_),
    .A2(_250_),
    .B(_237_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _630_ (.I(net87),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _631_ (.A1(net13),
    .A2(_234_),
    .ZN(_252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _632_ (.A1(_251_),
    .A2(_235_),
    .B(_252_),
    .C(_247_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _633_ (.I(net14),
    .Z(_253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _634_ (.A1(_253_),
    .A2(_230_),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _635_ (.A1(net88),
    .A2(_242_),
    .ZN(_255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _636_ (.A1(_254_),
    .A2(_255_),
    .B(_237_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _637_ (.I(net15),
    .Z(_256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _638_ (.A1(_256_),
    .A2(_229_),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _639_ (.A1(net89),
    .A2(_242_),
    .ZN(_258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _640_ (.I(net35),
    .Z(_259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _641_ (.I(_259_),
    .Z(_260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _642_ (.A1(_257_),
    .A2(_258_),
    .B(_260_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _643_ (.I(_210_),
    .Z(_261_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _644_ (.A1(_143_),
    .A2(_261_),
    .Z(_262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _645_ (.I(_262_),
    .Z(_263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _646_ (.A1(_226_),
    .A2(_263_),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _647_ (.A1(_143_),
    .A2(_211_),
    .ZN(_265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _648_ (.I(_265_),
    .Z(_266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _649_ (.A1(\DDRA[0] ),
    .A2(_266_),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _650_ (.A1(_264_),
    .A2(_267_),
    .B(_260_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _651_ (.I(net9),
    .Z(_268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _652_ (.A1(_268_),
    .A2(_263_),
    .ZN(_269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _653_ (.A1(\DDRA[1] ),
    .A2(_266_),
    .ZN(_270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _654_ (.A1(_269_),
    .A2(_270_),
    .B(_260_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _655_ (.A1(_240_),
    .A2(_263_),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _656_ (.A1(\DDRA[2] ),
    .A2(_266_),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _657_ (.A1(_271_),
    .A2(_272_),
    .B(_260_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _658_ (.I(net11),
    .Z(_273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _659_ (.A1(_273_),
    .A2(_263_),
    .ZN(_274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _660_ (.A1(\DDRA[3] ),
    .A2(_266_),
    .ZN(_275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _661_ (.I(_259_),
    .Z(_276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _662_ (.A1(_274_),
    .A2(_275_),
    .B(_276_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _663_ (.I(_262_),
    .Z(_277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _664_ (.A1(_248_),
    .A2(_277_),
    .ZN(_278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _665_ (.I(_265_),
    .Z(_279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _666_ (.A1(\DDRA[4] ),
    .A2(_279_),
    .ZN(_280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _667_ (.A1(_278_),
    .A2(_280_),
    .B(_276_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _668_ (.I(net13),
    .Z(_281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _669_ (.A1(_281_),
    .A2(_277_),
    .ZN(_282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _670_ (.A1(\DDRA[5] ),
    .A2(_279_),
    .ZN(_283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _671_ (.A1(_282_),
    .A2(_283_),
    .B(_276_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _672_ (.A1(_253_),
    .A2(_277_),
    .ZN(_284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _673_ (.A1(\DDRA[6] ),
    .A2(_279_),
    .ZN(_285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _674_ (.A1(_284_),
    .A2(_285_),
    .B(_276_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _675_ (.A1(_256_),
    .A2(_277_),
    .ZN(_286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _676_ (.A1(\DDRA[7] ),
    .A2(_279_),
    .ZN(_287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _677_ (.I(_259_),
    .Z(_288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _678_ (.A1(_286_),
    .A2(_287_),
    .B(_288_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _679_ (.A1(_135_),
    .A2(_116_),
    .A3(_118_),
    .A4(_132_),
    .ZN(_289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _680_ (.A1(_289_),
    .A2(_228_),
    .ZN(_290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _681_ (.I(_290_),
    .Z(_291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _682_ (.A1(_226_),
    .A2(_291_),
    .ZN(_292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _683_ (.A1(_127_),
    .A2(_210_),
    .ZN(_293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _684_ (.I(_293_),
    .Z(_294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _685_ (.A1(\DDRB[0] ),
    .A2(_294_),
    .ZN(_295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _686_ (.A1(_292_),
    .A2(_295_),
    .B(_288_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _687_ (.I(\DDRB[1] ),
    .ZN(_296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _688_ (.A1(net9),
    .A2(_293_),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _689_ (.A1(_296_),
    .A2(_294_),
    .B(_297_),
    .C(_247_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _690_ (.A1(_240_),
    .A2(_291_),
    .ZN(_298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _691_ (.A1(\DDRB[2] ),
    .A2(_294_),
    .ZN(_299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _692_ (.A1(_298_),
    .A2(_299_),
    .B(_288_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _693_ (.A1(_273_),
    .A2(_291_),
    .ZN(_300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _694_ (.A1(\DDRB[3] ),
    .A2(_294_),
    .ZN(_301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _695_ (.A1(_300_),
    .A2(_301_),
    .B(_288_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _696_ (.A1(_248_),
    .A2(_291_),
    .ZN(_302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _697_ (.I(_293_),
    .Z(_303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _698_ (.A1(\DDRB[4] ),
    .A2(_303_),
    .ZN(_304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _699_ (.I(_259_),
    .Z(_305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _700_ (.A1(_302_),
    .A2(_304_),
    .B(_305_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _701_ (.A1(_281_),
    .A2(_290_),
    .ZN(_306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _702_ (.A1(\DDRB[5] ),
    .A2(_303_),
    .ZN(_307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _703_ (.A1(_306_),
    .A2(_307_),
    .B(_305_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _704_ (.A1(_253_),
    .A2(_290_),
    .ZN(_308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _705_ (.A1(\DDRB[6] ),
    .A2(_303_),
    .ZN(_309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _706_ (.A1(_308_),
    .A2(_309_),
    .B(_305_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _707_ (.A1(_256_),
    .A2(_290_),
    .ZN(_310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _708_ (.A1(\DDRB[7] ),
    .A2(_303_),
    .ZN(_311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _709_ (.A1(_310_),
    .A2(_311_),
    .B(_305_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _710_ (.A1(_136_),
    .A2(_261_),
    .Z(_312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _711_ (.I(_312_),
    .Z(_313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _712_ (.A1(_226_),
    .A2(_313_),
    .ZN(_314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _713_ (.A1(_154_),
    .A2(_261_),
    .ZN(_315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _714_ (.I(_315_),
    .Z(_316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _715_ (.A1(\PORTA[0] ),
    .A2(_316_),
    .ZN(_317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _716_ (.I(net35),
    .Z(_318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _717_ (.I(_318_),
    .Z(_319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _718_ (.A1(_314_),
    .A2(_317_),
    .B(_319_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _719_ (.A1(_268_),
    .A2(_313_),
    .ZN(_320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _720_ (.A1(\PORTA[1] ),
    .A2(_316_),
    .ZN(_321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _721_ (.A1(_320_),
    .A2(_321_),
    .B(_319_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _722_ (.A1(_240_),
    .A2(_313_),
    .ZN(_322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _723_ (.A1(\PORTA[2] ),
    .A2(_316_),
    .ZN(_323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _724_ (.A1(_322_),
    .A2(_323_),
    .B(_319_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _725_ (.A1(_273_),
    .A2(_313_),
    .ZN(_324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _726_ (.A1(\PORTA[3] ),
    .A2(_316_),
    .ZN(_325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _727_ (.A1(_324_),
    .A2(_325_),
    .B(_319_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _728_ (.I(_312_),
    .Z(_326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _729_ (.A1(_248_),
    .A2(_326_),
    .ZN(_327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _730_ (.I(_315_),
    .Z(_328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _731_ (.A1(\PORTA[4] ),
    .A2(_328_),
    .ZN(_329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _732_ (.I(_318_),
    .Z(_330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _733_ (.A1(_327_),
    .A2(_329_),
    .B(_330_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _734_ (.A1(_281_),
    .A2(_326_),
    .ZN(_331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _735_ (.A1(\PORTA[5] ),
    .A2(_328_),
    .ZN(_332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _736_ (.A1(_331_),
    .A2(_332_),
    .B(_330_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _737_ (.A1(_253_),
    .A2(_326_),
    .ZN(_333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _738_ (.A1(\PORTA[6] ),
    .A2(_328_),
    .ZN(_334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _739_ (.A1(_333_),
    .A2(_334_),
    .B(_330_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _740_ (.A1(_256_),
    .A2(_326_),
    .ZN(_335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _741_ (.A1(\PORTA[7] ),
    .A2(_328_),
    .ZN(_336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _742_ (.A1(_335_),
    .A2(_336_),
    .B(_330_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _743_ (.A1(_129_),
    .A2(_232_),
    .Z(_337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _744_ (.I(_337_),
    .Z(_338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _745_ (.A1(_208_),
    .A2(_338_),
    .ZN(_339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _746_ (.A1(_129_),
    .A2(_261_),
    .ZN(_340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _747_ (.I(_340_),
    .Z(_341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _748_ (.A1(\PORTB[0] ),
    .A2(_341_),
    .ZN(_342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _749_ (.I(_318_),
    .Z(_343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _750_ (.A1(_339_),
    .A2(_342_),
    .B(_343_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _751_ (.A1(_268_),
    .A2(_338_),
    .ZN(_344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _752_ (.A1(\PORTB[1] ),
    .A2(_341_),
    .ZN(_345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _753_ (.A1(_344_),
    .A2(_345_),
    .B(_343_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _754_ (.A1(net10),
    .A2(_338_),
    .ZN(_346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _755_ (.A1(\PORTB[2] ),
    .A2(_341_),
    .ZN(_347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _756_ (.A1(_346_),
    .A2(_347_),
    .B(_343_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _757_ (.A1(_273_),
    .A2(_338_),
    .ZN(_348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _758_ (.A1(\PORTB[3] ),
    .A2(_341_),
    .ZN(_349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _759_ (.A1(_348_),
    .A2(_349_),
    .B(_343_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _760_ (.I(_337_),
    .Z(_350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _761_ (.A1(net12),
    .A2(_350_),
    .ZN(_351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _762_ (.I(_340_),
    .Z(_352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _763_ (.A1(\PORTB[4] ),
    .A2(_352_),
    .ZN(_353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _764_ (.I(_318_),
    .Z(_354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _765_ (.A1(_351_),
    .A2(_353_),
    .B(_354_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _766_ (.A1(_281_),
    .A2(_350_),
    .ZN(_355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _767_ (.A1(\PORTB[5] ),
    .A2(_352_),
    .ZN(_356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _768_ (.A1(_355_),
    .A2(_356_),
    .B(_354_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _769_ (.A1(_216_),
    .A2(_350_),
    .ZN(_357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _770_ (.A1(\PORTB[6] ),
    .A2(_352_),
    .ZN(_358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _771_ (.A1(_357_),
    .A2(_358_),
    .B(_354_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _772_ (.A1(_222_),
    .A2(_350_),
    .ZN(_359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _773_ (.A1(\PORTB[7] ),
    .A2(_352_),
    .ZN(_360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _774_ (.A1(_359_),
    .A2(_360_),
    .B(_354_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _775_ (.A1(_138_),
    .A2(_210_),
    .ZN(_361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _776_ (.I(_361_),
    .Z(_362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _777_ (.I(_362_),
    .Z(_363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _778_ (.A1(_208_),
    .A2(_362_),
    .ZN(_364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _779_ (.A1(_070_),
    .A2(_363_),
    .B(_364_),
    .C(_247_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _780_ (.A1(_138_),
    .A2(_232_),
    .Z(_365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _781_ (.I(_365_),
    .Z(_366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _782_ (.A1(_268_),
    .A2(_366_),
    .ZN(_367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _783_ (.A1(\SPA[1] ),
    .A2(_363_),
    .ZN(_368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _784_ (.I(_246_),
    .Z(_369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _785_ (.A1(_367_),
    .A2(_368_),
    .B(_369_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _786_ (.A1(net10),
    .A2(_362_),
    .ZN(_370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _787_ (.I(_246_),
    .Z(_371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _788_ (.A1(_073_),
    .A2(_363_),
    .B(_370_),
    .C(_371_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _789_ (.A1(net11),
    .A2(_366_),
    .ZN(_372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _790_ (.I(_361_),
    .Z(_373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _791_ (.A1(\SPA[3] ),
    .A2(_373_),
    .ZN(_374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _792_ (.A1(_372_),
    .A2(_374_),
    .B(_369_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _793_ (.A1(net12),
    .A2(_366_),
    .ZN(_375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _794_ (.A1(\SPA[4] ),
    .A2(_373_),
    .ZN(_376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _795_ (.A1(_375_),
    .A2(_376_),
    .B(_369_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _796_ (.A1(net13),
    .A2(_366_),
    .ZN(_377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _797_ (.A1(\SPA[5] ),
    .A2(_373_),
    .ZN(_378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _798_ (.A1(_377_),
    .A2(_378_),
    .B(_369_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _799_ (.A1(_216_),
    .A2(_365_),
    .ZN(_379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _800_ (.A1(\SPA[6] ),
    .A2(_373_),
    .ZN(_380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _801_ (.A1(_379_),
    .A2(_380_),
    .B(_101_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _802_ (.A1(_222_),
    .A2(_362_),
    .ZN(_381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _803_ (.A1(_079_),
    .A2(_363_),
    .B(_381_),
    .C(_371_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _804_ (.A1(_111_),
    .A2(_232_),
    .ZN(_382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _805_ (.I(_382_),
    .Z(_383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _806_ (.I(_382_),
    .Z(_384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _807_ (.A1(_208_),
    .A2(_384_),
    .ZN(_385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _808_ (.A1(_082_),
    .A2(_383_),
    .B(_385_),
    .C(_371_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _809_ (.I(\SPB[1] ),
    .ZN(_386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _810_ (.A1(net9),
    .A2(_384_),
    .ZN(_387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _811_ (.A1(_386_),
    .A2(_383_),
    .B(_387_),
    .C(_371_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _812_ (.A1(net10),
    .A2(_384_),
    .ZN(_388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _813_ (.I(_246_),
    .Z(_389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _814_ (.A1(_085_),
    .A2(_383_),
    .B(_388_),
    .C(_389_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _815_ (.A1(net11),
    .A2(_384_),
    .ZN(_390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _816_ (.A1(_087_),
    .A2(_383_),
    .B(_390_),
    .C(_389_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _817_ (.I(_382_),
    .Z(_391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _818_ (.I(_382_),
    .Z(_392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _819_ (.A1(net12),
    .A2(_392_),
    .ZN(_393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _820_ (.A1(_089_),
    .A2(_391_),
    .B(_393_),
    .C(_389_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _821_ (.A1(net13),
    .A2(_392_),
    .ZN(_394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _822_ (.A1(_091_),
    .A2(_391_),
    .B(_394_),
    .C(_389_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _823_ (.A1(_216_),
    .A2(_392_),
    .ZN(_395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _824_ (.A1(_093_),
    .A2(_391_),
    .B(_395_),
    .C(_148_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _825_ (.A1(_222_),
    .A2(_392_),
    .ZN(_396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _826_ (.A1(_095_),
    .A2(_391_),
    .B(_396_),
    .C(_148_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _827_ (.A1(_221_),
    .A2(_213_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _828_ (.A1(_221_),
    .A2(_218_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _829_ (.D(_000_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(last_irq7_trigger));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _830_ (.D(_001_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _831_ (.D(_002_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _832_ (.D(_003_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _833_ (.D(_004_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _834_ (.D(_005_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _835_ (.D(_006_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _836_ (.D(_007_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _837_ (.D(_008_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net46));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _838_ (.D(_009_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(net79));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _839_ (.D(_010_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net80));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _840_ (.D(_011_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(net81));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _841_ (.D(_012_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net82));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _842_ (.D(_013_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net83));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _843_ (.D(_014_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net84));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _844_ (.D(_015_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net85));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _845_ (.D(_016_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net86));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _846_ (.D(_017_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net87));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _847_ (.D(_018_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net88));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _848_ (.D(_019_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net89));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _849_ (.D(_020_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _850_ (.D(_021_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _851_ (.D(_022_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _852_ (.D(_023_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _853_ (.D(_024_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _854_ (.D(_025_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _855_ (.D(_026_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _856_ (.D(_027_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _857_ (.D(_028_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _858_ (.D(_029_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _859_ (.D(_030_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _860_ (.D(_031_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _861_ (.D(_032_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _862_ (.D(_033_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\DDRB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _863_ (.D(_034_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\DDRB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _864_ (.D(_035_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\DDRB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _865_ (.D(_036_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\PORTA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _866_ (.D(_037_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\PORTA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _867_ (.D(_038_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\PORTA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _868_ (.D(_039_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\PORTA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _869_ (.D(_040_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _870_ (.D(_041_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _871_ (.D(_042_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _872_ (.D(_043_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _873_ (.D(_044_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _874_ (.D(_045_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _875_ (.D(_046_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _876_ (.D(_047_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _877_ (.D(_048_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _878_ (.D(_049_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _879_ (.D(_050_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _880_ (.D(_051_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _881_ (.D(_052_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(\SPA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _882_ (.D(_053_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\SPA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _883_ (.D(_054_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\SPA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _884_ (.D(_055_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\SPA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _885_ (.D(_056_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\SPA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _886_ (.D(_057_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\SPA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _887_ (.D(_058_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\SPA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _888_ (.D(_059_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _889_ (.D(_060_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _890_ (.D(_061_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _891_ (.D(_062_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _892_ (.D(_063_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _893_ (.D(_064_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\SPB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _894_ (.D(_065_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _895_ (.D(_066_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\SPB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _896_ (.D(_067_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\SPB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _897_ (.D(_068_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(last_irq0_trigger));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _898_ (.D(_069_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(last_irg6_trigger));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold1 (.I(net88),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold2 (.I(net85),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold3 (.I(net83),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold4 (.I(net82),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold5 (.I(net86),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold6 (.I(net87),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold7 (.I(net84),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold8 (.I(net89),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(TXD),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input10 (.I(data_in[2]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input11 (.I(data_in[3]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input12 (.I(data_in[4]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input13 (.I(data_in[5]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(data_in[6]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(data_in[7]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input16 (.I(io_in[0]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(io_in[10]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(io_in[11]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(io_in[12]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input2 (.I(addr[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(io_in[13]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(io_in[14]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(io_in[15]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(io_in[1]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(io_in[2]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(io_in[3]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(io_in[4]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(io_in[5]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(io_in[6]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input29 (.I(io_in[7]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(addr[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(io_in[8]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(io_in[9]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(pwm0),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(pwm1),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(pwm2),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input35 (.I(rst),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input36 (.I(tmr0_o),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(tmr1_o),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(addr[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(addr[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input6 (.I(bus_cyc),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(bus_we),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(data_in[0]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input9 (.I(data_in[1]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output38 (.I(net38),
    .Z(RXD));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output39 (.I(net39),
    .Z(data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output40 (.I(net40),
    .Z(data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output41 (.I(net41),
    .Z(data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output42 (.I(net42),
    .Z(data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output43 (.I(net43),
    .Z(data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output44 (.I(net44),
    .Z(data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output45 (.I(net45),
    .Z(data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output46 (.I(net46),
    .Z(data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output47 (.I(net47),
    .Z(io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output48 (.I(net48),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output49 (.I(net49),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output50 (.I(net50),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output51 (.I(net51),
    .Z(io_oeb[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output52 (.I(net52),
    .Z(io_oeb[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output53 (.I(net53),
    .Z(io_oeb[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output54 (.I(net54),
    .Z(io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output55 (.I(net55),
    .Z(io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output56 (.I(net56),
    .Z(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output57 (.I(net57),
    .Z(io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output58 (.I(net58),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output59 (.I(net59),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output60 (.I(net60),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output61 (.I(net61),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output62 (.I(net62),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output63 (.I(net63),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output64 (.I(net64),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output65 (.I(net65),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output66 (.I(net66),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output67 (.I(net67),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output68 (.I(net68),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output69 (.I(net69),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output70 (.I(net70),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output71 (.I(net71),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output72 (.I(net72),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output73 (.I(net73),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output74 (.I(net74),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output75 (.I(net75),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output76 (.I(net76),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output77 (.I(net77),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output78 (.I(net78),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output79 (.I(net79),
    .Z(irq0));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output80 (.I(net80),
    .Z(irq6));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output81 (.I(net81),
    .Z(irq7));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output82 (.I(net95),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output83 (.I(net94),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output84 (.I(net98),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output85 (.I(net93),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output86 (.I(net96),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output87 (.I(net97),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output88 (.I(net92),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output89 (.I(net99),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output90 (.I(net90),
    .Z(tmr0_clk));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output91 (.I(net91),
    .Z(tmr1_clk));
endmodule

