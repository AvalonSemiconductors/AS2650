// This is the unpowered netlist.
module sid_top (DAC_clk,
    DAC_dat_1,
    DAC_dat_2,
    DAC_le,
    bus_cyc,
    bus_we,
    clk,
    rst,
    addr,
    bus_in,
    bus_out);
 output DAC_clk;
 output DAC_dat_1;
 output DAC_dat_2;
 output DAC_le;
 input bus_cyc;
 input bus_we;
 input clk;
 input rst;
 input [4:0] addr;
 input [7:0] bus_in;
 output [7:0] bus_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire \channels.accum[0][0] ;
 wire \channels.accum[0][10] ;
 wire \channels.accum[0][11] ;
 wire \channels.accum[0][12] ;
 wire \channels.accum[0][13] ;
 wire \channels.accum[0][14] ;
 wire \channels.accum[0][15] ;
 wire \channels.accum[0][16] ;
 wire \channels.accum[0][17] ;
 wire \channels.accum[0][18] ;
 wire \channels.accum[0][19] ;
 wire \channels.accum[0][1] ;
 wire \channels.accum[0][20] ;
 wire \channels.accum[0][21] ;
 wire \channels.accum[0][22] ;
 wire \channels.accum[0][23] ;
 wire \channels.accum[0][2] ;
 wire \channels.accum[0][3] ;
 wire \channels.accum[0][4] ;
 wire \channels.accum[0][5] ;
 wire \channels.accum[0][6] ;
 wire \channels.accum[0][7] ;
 wire \channels.accum[0][8] ;
 wire \channels.accum[0][9] ;
 wire \channels.accum[1][0] ;
 wire \channels.accum[1][10] ;
 wire \channels.accum[1][11] ;
 wire \channels.accum[1][12] ;
 wire \channels.accum[1][13] ;
 wire \channels.accum[1][14] ;
 wire \channels.accum[1][15] ;
 wire \channels.accum[1][16] ;
 wire \channels.accum[1][17] ;
 wire \channels.accum[1][18] ;
 wire \channels.accum[1][19] ;
 wire \channels.accum[1][1] ;
 wire \channels.accum[1][20] ;
 wire \channels.accum[1][21] ;
 wire \channels.accum[1][22] ;
 wire \channels.accum[1][23] ;
 wire \channels.accum[1][2] ;
 wire \channels.accum[1][3] ;
 wire \channels.accum[1][4] ;
 wire \channels.accum[1][5] ;
 wire \channels.accum[1][6] ;
 wire \channels.accum[1][7] ;
 wire \channels.accum[1][8] ;
 wire \channels.accum[1][9] ;
 wire \channels.accum[2][0] ;
 wire \channels.accum[2][10] ;
 wire \channels.accum[2][11] ;
 wire \channels.accum[2][12] ;
 wire \channels.accum[2][13] ;
 wire \channels.accum[2][14] ;
 wire \channels.accum[2][15] ;
 wire \channels.accum[2][16] ;
 wire \channels.accum[2][17] ;
 wire \channels.accum[2][18] ;
 wire \channels.accum[2][19] ;
 wire \channels.accum[2][1] ;
 wire \channels.accum[2][20] ;
 wire \channels.accum[2][21] ;
 wire \channels.accum[2][22] ;
 wire \channels.accum[2][23] ;
 wire \channels.accum[2][2] ;
 wire \channels.accum[2][3] ;
 wire \channels.accum[2][4] ;
 wire \channels.accum[2][5] ;
 wire \channels.accum[2][6] ;
 wire \channels.accum[2][7] ;
 wire \channels.accum[2][8] ;
 wire \channels.accum[2][9] ;
 wire \channels.accum[3][0] ;
 wire \channels.accum[3][10] ;
 wire \channels.accum[3][11] ;
 wire \channels.accum[3][12] ;
 wire \channels.accum[3][13] ;
 wire \channels.accum[3][14] ;
 wire \channels.accum[3][15] ;
 wire \channels.accum[3][16] ;
 wire \channels.accum[3][17] ;
 wire \channels.accum[3][18] ;
 wire \channels.accum[3][19] ;
 wire \channels.accum[3][1] ;
 wire \channels.accum[3][20] ;
 wire \channels.accum[3][21] ;
 wire \channels.accum[3][22] ;
 wire \channels.accum[3][23] ;
 wire \channels.accum[3][2] ;
 wire \channels.accum[3][3] ;
 wire \channels.accum[3][4] ;
 wire \channels.accum[3][5] ;
 wire \channels.accum[3][6] ;
 wire \channels.accum[3][7] ;
 wire \channels.accum[3][8] ;
 wire \channels.accum[3][9] ;
 wire \channels.adsr_state[0][0] ;
 wire \channels.adsr_state[0][1] ;
 wire \channels.adsr_state[1][0] ;
 wire \channels.adsr_state[1][1] ;
 wire \channels.adsr_state[2][0] ;
 wire \channels.adsr_state[2][1] ;
 wire \channels.adsr_state[3][0] ;
 wire \channels.adsr_state[3][1] ;
 wire \channels.atk_dec1[0] ;
 wire \channels.atk_dec1[1] ;
 wire \channels.atk_dec1[2] ;
 wire \channels.atk_dec1[3] ;
 wire \channels.atk_dec1[4] ;
 wire \channels.atk_dec1[5] ;
 wire \channels.atk_dec1[6] ;
 wire \channels.atk_dec1[7] ;
 wire \channels.atk_dec2[0] ;
 wire \channels.atk_dec2[1] ;
 wire \channels.atk_dec2[2] ;
 wire \channels.atk_dec2[3] ;
 wire \channels.atk_dec2[4] ;
 wire \channels.atk_dec2[5] ;
 wire \channels.atk_dec2[6] ;
 wire \channels.atk_dec2[7] ;
 wire \channels.atk_dec3[0] ;
 wire \channels.atk_dec3[1] ;
 wire \channels.atk_dec3[2] ;
 wire \channels.atk_dec3[3] ;
 wire \channels.atk_dec3[4] ;
 wire \channels.atk_dec3[5] ;
 wire \channels.atk_dec3[6] ;
 wire \channels.atk_dec3[7] ;
 wire \channels.ch3_env[0] ;
 wire \channels.ch3_env[1] ;
 wire \channels.ch3_env[2] ;
 wire \channels.ch3_env[3] ;
 wire \channels.ch3_env[4] ;
 wire \channels.ch3_env[5] ;
 wire \channels.ch3_env[6] ;
 wire \channels.ch3_env[7] ;
 wire \channels.clk_div[0] ;
 wire \channels.clk_div[1] ;
 wire \channels.clk_div[2] ;
 wire \channels.ctrl_reg1[0] ;
 wire \channels.ctrl_reg1[1] ;
 wire \channels.ctrl_reg1[2] ;
 wire \channels.ctrl_reg1[3] ;
 wire \channels.ctrl_reg1[4] ;
 wire \channels.ctrl_reg1[5] ;
 wire \channels.ctrl_reg1[6] ;
 wire \channels.ctrl_reg1[7] ;
 wire \channels.ctrl_reg2[0] ;
 wire \channels.ctrl_reg2[1] ;
 wire \channels.ctrl_reg2[2] ;
 wire \channels.ctrl_reg2[3] ;
 wire \channels.ctrl_reg2[4] ;
 wire \channels.ctrl_reg2[5] ;
 wire \channels.ctrl_reg2[6] ;
 wire \channels.ctrl_reg2[7] ;
 wire \channels.ctrl_reg3[0] ;
 wire \channels.ctrl_reg3[1] ;
 wire \channels.ctrl_reg3[2] ;
 wire \channels.ctrl_reg3[3] ;
 wire \channels.ctrl_reg3[4] ;
 wire \channels.ctrl_reg3[5] ;
 wire \channels.ctrl_reg3[6] ;
 wire \channels.ctrl_reg3[7] ;
 wire \channels.env_counter[0][0] ;
 wire \channels.env_counter[0][10] ;
 wire \channels.env_counter[0][11] ;
 wire \channels.env_counter[0][12] ;
 wire \channels.env_counter[0][13] ;
 wire \channels.env_counter[0][14] ;
 wire \channels.env_counter[0][1] ;
 wire \channels.env_counter[0][2] ;
 wire \channels.env_counter[0][3] ;
 wire \channels.env_counter[0][4] ;
 wire \channels.env_counter[0][5] ;
 wire \channels.env_counter[0][6] ;
 wire \channels.env_counter[0][7] ;
 wire \channels.env_counter[0][8] ;
 wire \channels.env_counter[0][9] ;
 wire \channels.env_counter[1][0] ;
 wire \channels.env_counter[1][10] ;
 wire \channels.env_counter[1][11] ;
 wire \channels.env_counter[1][12] ;
 wire \channels.env_counter[1][13] ;
 wire \channels.env_counter[1][14] ;
 wire \channels.env_counter[1][1] ;
 wire \channels.env_counter[1][2] ;
 wire \channels.env_counter[1][3] ;
 wire \channels.env_counter[1][4] ;
 wire \channels.env_counter[1][5] ;
 wire \channels.env_counter[1][6] ;
 wire \channels.env_counter[1][7] ;
 wire \channels.env_counter[1][8] ;
 wire \channels.env_counter[1][9] ;
 wire \channels.env_counter[2][0] ;
 wire \channels.env_counter[2][10] ;
 wire \channels.env_counter[2][11] ;
 wire \channels.env_counter[2][12] ;
 wire \channels.env_counter[2][13] ;
 wire \channels.env_counter[2][14] ;
 wire \channels.env_counter[2][1] ;
 wire \channels.env_counter[2][2] ;
 wire \channels.env_counter[2][3] ;
 wire \channels.env_counter[2][4] ;
 wire \channels.env_counter[2][5] ;
 wire \channels.env_counter[2][6] ;
 wire \channels.env_counter[2][7] ;
 wire \channels.env_counter[2][8] ;
 wire \channels.env_counter[2][9] ;
 wire \channels.env_counter[3][0] ;
 wire \channels.env_counter[3][10] ;
 wire \channels.env_counter[3][11] ;
 wire \channels.env_counter[3][12] ;
 wire \channels.env_counter[3][13] ;
 wire \channels.env_counter[3][14] ;
 wire \channels.env_counter[3][1] ;
 wire \channels.env_counter[3][2] ;
 wire \channels.env_counter[3][3] ;
 wire \channels.env_counter[3][4] ;
 wire \channels.env_counter[3][5] ;
 wire \channels.env_counter[3][6] ;
 wire \channels.env_counter[3][7] ;
 wire \channels.env_counter[3][8] ;
 wire \channels.env_counter[3][9] ;
 wire \channels.env_vol[0][0] ;
 wire \channels.env_vol[0][1] ;
 wire \channels.env_vol[0][2] ;
 wire \channels.env_vol[0][3] ;
 wire \channels.env_vol[0][4] ;
 wire \channels.env_vol[0][5] ;
 wire \channels.env_vol[0][6] ;
 wire \channels.env_vol[0][7] ;
 wire \channels.env_vol[1][0] ;
 wire \channels.env_vol[1][1] ;
 wire \channels.env_vol[1][2] ;
 wire \channels.env_vol[1][3] ;
 wire \channels.env_vol[1][4] ;
 wire \channels.env_vol[1][5] ;
 wire \channels.env_vol[1][6] ;
 wire \channels.env_vol[1][7] ;
 wire \channels.env_vol[3][0] ;
 wire \channels.env_vol[3][1] ;
 wire \channels.env_vol[3][2] ;
 wire \channels.env_vol[3][3] ;
 wire \channels.env_vol[3][4] ;
 wire \channels.env_vol[3][5] ;
 wire \channels.env_vol[3][6] ;
 wire \channels.env_vol[3][7] ;
 wire \channels.exp_counter[0][0] ;
 wire \channels.exp_counter[0][1] ;
 wire \channels.exp_counter[0][2] ;
 wire \channels.exp_counter[0][3] ;
 wire \channels.exp_counter[0][4] ;
 wire \channels.exp_counter[1][0] ;
 wire \channels.exp_counter[1][1] ;
 wire \channels.exp_counter[1][2] ;
 wire \channels.exp_counter[1][3] ;
 wire \channels.exp_counter[1][4] ;
 wire \channels.exp_counter[2][0] ;
 wire \channels.exp_counter[2][1] ;
 wire \channels.exp_counter[2][2] ;
 wire \channels.exp_counter[2][3] ;
 wire \channels.exp_counter[2][4] ;
 wire \channels.exp_counter[3][0] ;
 wire \channels.exp_counter[3][1] ;
 wire \channels.exp_counter[3][2] ;
 wire \channels.exp_counter[3][3] ;
 wire \channels.exp_counter[3][4] ;
 wire \channels.exp_periods[0][0] ;
 wire \channels.exp_periods[0][1] ;
 wire \channels.exp_periods[0][2] ;
 wire \channels.exp_periods[0][3] ;
 wire \channels.exp_periods[0][4] ;
 wire \channels.exp_periods[1][0] ;
 wire \channels.exp_periods[1][1] ;
 wire \channels.exp_periods[1][2] ;
 wire \channels.exp_periods[1][3] ;
 wire \channels.exp_periods[1][4] ;
 wire \channels.exp_periods[2][0] ;
 wire \channels.exp_periods[2][1] ;
 wire \channels.exp_periods[2][2] ;
 wire \channels.exp_periods[2][3] ;
 wire \channels.exp_periods[2][4] ;
 wire \channels.exp_periods[3][0] ;
 wire \channels.exp_periods[3][1] ;
 wire \channels.exp_periods[3][2] ;
 wire \channels.exp_periods[3][3] ;
 wire \channels.exp_periods[3][4] ;
 wire \channels.freq1[0] ;
 wire \channels.freq1[10] ;
 wire \channels.freq1[11] ;
 wire \channels.freq1[12] ;
 wire \channels.freq1[13] ;
 wire \channels.freq1[14] ;
 wire \channels.freq1[15] ;
 wire \channels.freq1[1] ;
 wire \channels.freq1[2] ;
 wire \channels.freq1[3] ;
 wire \channels.freq1[4] ;
 wire \channels.freq1[5] ;
 wire \channels.freq1[6] ;
 wire \channels.freq1[7] ;
 wire \channels.freq1[8] ;
 wire \channels.freq1[9] ;
 wire \channels.freq2[0] ;
 wire \channels.freq2[10] ;
 wire \channels.freq2[11] ;
 wire \channels.freq2[12] ;
 wire \channels.freq2[13] ;
 wire \channels.freq2[14] ;
 wire \channels.freq2[15] ;
 wire \channels.freq2[1] ;
 wire \channels.freq2[2] ;
 wire \channels.freq2[3] ;
 wire \channels.freq2[4] ;
 wire \channels.freq2[5] ;
 wire \channels.freq2[6] ;
 wire \channels.freq2[7] ;
 wire \channels.freq2[8] ;
 wire \channels.freq2[9] ;
 wire \channels.freq3[0] ;
 wire \channels.freq3[10] ;
 wire \channels.freq3[11] ;
 wire \channels.freq3[12] ;
 wire \channels.freq3[13] ;
 wire \channels.freq3[14] ;
 wire \channels.freq3[15] ;
 wire \channels.freq3[1] ;
 wire \channels.freq3[2] ;
 wire \channels.freq3[3] ;
 wire \channels.freq3[4] ;
 wire \channels.freq3[5] ;
 wire \channels.freq3[6] ;
 wire \channels.freq3[7] ;
 wire \channels.freq3[8] ;
 wire \channels.freq3[9] ;
 wire \channels.lfsr[0][0] ;
 wire \channels.lfsr[0][10] ;
 wire \channels.lfsr[0][11] ;
 wire \channels.lfsr[0][12] ;
 wire \channels.lfsr[0][13] ;
 wire \channels.lfsr[0][14] ;
 wire \channels.lfsr[0][15] ;
 wire \channels.lfsr[0][16] ;
 wire \channels.lfsr[0][17] ;
 wire \channels.lfsr[0][18] ;
 wire \channels.lfsr[0][19] ;
 wire \channels.lfsr[0][1] ;
 wire \channels.lfsr[0][20] ;
 wire \channels.lfsr[0][21] ;
 wire \channels.lfsr[0][22] ;
 wire \channels.lfsr[0][2] ;
 wire \channels.lfsr[0][3] ;
 wire \channels.lfsr[0][4] ;
 wire \channels.lfsr[0][5] ;
 wire \channels.lfsr[0][6] ;
 wire \channels.lfsr[0][7] ;
 wire \channels.lfsr[0][8] ;
 wire \channels.lfsr[0][9] ;
 wire \channels.lfsr[1][0] ;
 wire \channels.lfsr[1][10] ;
 wire \channels.lfsr[1][11] ;
 wire \channels.lfsr[1][12] ;
 wire \channels.lfsr[1][13] ;
 wire \channels.lfsr[1][14] ;
 wire \channels.lfsr[1][15] ;
 wire \channels.lfsr[1][16] ;
 wire \channels.lfsr[1][17] ;
 wire \channels.lfsr[1][18] ;
 wire \channels.lfsr[1][19] ;
 wire \channels.lfsr[1][1] ;
 wire \channels.lfsr[1][20] ;
 wire \channels.lfsr[1][21] ;
 wire \channels.lfsr[1][22] ;
 wire \channels.lfsr[1][2] ;
 wire \channels.lfsr[1][3] ;
 wire \channels.lfsr[1][4] ;
 wire \channels.lfsr[1][5] ;
 wire \channels.lfsr[1][6] ;
 wire \channels.lfsr[1][7] ;
 wire \channels.lfsr[1][8] ;
 wire \channels.lfsr[1][9] ;
 wire \channels.lfsr[2][0] ;
 wire \channels.lfsr[2][10] ;
 wire \channels.lfsr[2][11] ;
 wire \channels.lfsr[2][12] ;
 wire \channels.lfsr[2][13] ;
 wire \channels.lfsr[2][14] ;
 wire \channels.lfsr[2][15] ;
 wire \channels.lfsr[2][16] ;
 wire \channels.lfsr[2][17] ;
 wire \channels.lfsr[2][18] ;
 wire \channels.lfsr[2][19] ;
 wire \channels.lfsr[2][1] ;
 wire \channels.lfsr[2][20] ;
 wire \channels.lfsr[2][21] ;
 wire \channels.lfsr[2][22] ;
 wire \channels.lfsr[2][2] ;
 wire \channels.lfsr[2][3] ;
 wire \channels.lfsr[2][4] ;
 wire \channels.lfsr[2][5] ;
 wire \channels.lfsr[2][6] ;
 wire \channels.lfsr[2][7] ;
 wire \channels.lfsr[2][8] ;
 wire \channels.lfsr[2][9] ;
 wire \channels.lfsr[3][0] ;
 wire \channels.lfsr[3][10] ;
 wire \channels.lfsr[3][11] ;
 wire \channels.lfsr[3][12] ;
 wire \channels.lfsr[3][13] ;
 wire \channels.lfsr[3][14] ;
 wire \channels.lfsr[3][15] ;
 wire \channels.lfsr[3][16] ;
 wire \channels.lfsr[3][17] ;
 wire \channels.lfsr[3][18] ;
 wire \channels.lfsr[3][19] ;
 wire \channels.lfsr[3][1] ;
 wire \channels.lfsr[3][20] ;
 wire \channels.lfsr[3][21] ;
 wire \channels.lfsr[3][22] ;
 wire \channels.lfsr[3][2] ;
 wire \channels.lfsr[3][3] ;
 wire \channels.lfsr[3][4] ;
 wire \channels.lfsr[3][5] ;
 wire \channels.lfsr[3][6] ;
 wire \channels.lfsr[3][7] ;
 wire \channels.lfsr[3][8] ;
 wire \channels.lfsr[3][9] ;
 wire \channels.pw1[0] ;
 wire \channels.pw1[10] ;
 wire \channels.pw1[11] ;
 wire \channels.pw1[1] ;
 wire \channels.pw1[2] ;
 wire \channels.pw1[3] ;
 wire \channels.pw1[4] ;
 wire \channels.pw1[5] ;
 wire \channels.pw1[6] ;
 wire \channels.pw1[7] ;
 wire \channels.pw1[8] ;
 wire \channels.pw1[9] ;
 wire \channels.pw2[0] ;
 wire \channels.pw2[10] ;
 wire \channels.pw2[11] ;
 wire \channels.pw2[1] ;
 wire \channels.pw2[2] ;
 wire \channels.pw2[3] ;
 wire \channels.pw2[4] ;
 wire \channels.pw2[5] ;
 wire \channels.pw2[6] ;
 wire \channels.pw2[7] ;
 wire \channels.pw2[8] ;
 wire \channels.pw2[9] ;
 wire \channels.pw3[0] ;
 wire \channels.pw3[10] ;
 wire \channels.pw3[11] ;
 wire \channels.pw3[1] ;
 wire \channels.pw3[2] ;
 wire \channels.pw3[3] ;
 wire \channels.pw3[4] ;
 wire \channels.pw3[5] ;
 wire \channels.pw3[6] ;
 wire \channels.pw3[7] ;
 wire \channels.pw3[8] ;
 wire \channels.pw3[9] ;
 wire \channels.ring_outs[0] ;
 wire \channels.ring_outs[1] ;
 wire \channels.ring_outs[2] ;
 wire \channels.sample1[0] ;
 wire \channels.sample1[10] ;
 wire \channels.sample1[11] ;
 wire \channels.sample1[1] ;
 wire \channels.sample1[2] ;
 wire \channels.sample1[3] ;
 wire \channels.sample1[4] ;
 wire \channels.sample1[5] ;
 wire \channels.sample1[6] ;
 wire \channels.sample1[7] ;
 wire \channels.sample1[8] ;
 wire \channels.sample1[9] ;
 wire \channels.sample2[0] ;
 wire \channels.sample2[10] ;
 wire \channels.sample2[11] ;
 wire \channels.sample2[1] ;
 wire \channels.sample2[2] ;
 wire \channels.sample2[3] ;
 wire \channels.sample2[4] ;
 wire \channels.sample2[5] ;
 wire \channels.sample2[6] ;
 wire \channels.sample2[7] ;
 wire \channels.sample2[8] ;
 wire \channels.sample2[9] ;
 wire \channels.sample3[0] ;
 wire \channels.sample3[10] ;
 wire \channels.sample3[11] ;
 wire \channels.sample3[1] ;
 wire \channels.sample3[2] ;
 wire \channels.sample3[3] ;
 wire \channels.sample3[4] ;
 wire \channels.sample3[5] ;
 wire \channels.sample3[6] ;
 wire \channels.sample3[7] ;
 wire \channels.sample3[8] ;
 wire \channels.sample3[9] ;
 wire \channels.sus_rel1[0] ;
 wire \channels.sus_rel1[1] ;
 wire \channels.sus_rel1[2] ;
 wire \channels.sus_rel1[3] ;
 wire \channels.sus_rel1[4] ;
 wire \channels.sus_rel1[5] ;
 wire \channels.sus_rel1[6] ;
 wire \channels.sus_rel1[7] ;
 wire \channels.sus_rel2[0] ;
 wire \channels.sus_rel2[1] ;
 wire \channels.sus_rel2[2] ;
 wire \channels.sus_rel2[3] ;
 wire \channels.sus_rel2[4] ;
 wire \channels.sus_rel2[5] ;
 wire \channels.sus_rel2[6] ;
 wire \channels.sus_rel2[7] ;
 wire \channels.sus_rel3[0] ;
 wire \channels.sus_rel3[1] ;
 wire \channels.sus_rel3[2] ;
 wire \channels.sus_rel3[3] ;
 wire \channels.sus_rel3[4] ;
 wire \channels.sus_rel3[5] ;
 wire \channels.sus_rel3[6] ;
 wire \channels.sus_rel3[7] ;
 wire \channels.sync_outs[0] ;
 wire \channels.sync_outs[1] ;
 wire \channels.sync_outs[2] ;
 wire \clk_ctr[0] ;
 wire \clk_ctr[1] ;
 wire \clk_trg[0] ;
 wire \clk_trg[1] ;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_9_clk;
 wire \filters.band[0] ;
 wire \filters.band[10] ;
 wire \filters.band[11] ;
 wire \filters.band[12] ;
 wire \filters.band[13] ;
 wire \filters.band[14] ;
 wire \filters.band[15] ;
 wire \filters.band[16] ;
 wire \filters.band[17] ;
 wire \filters.band[18] ;
 wire \filters.band[19] ;
 wire \filters.band[1] ;
 wire \filters.band[20] ;
 wire \filters.band[21] ;
 wire \filters.band[22] ;
 wire \filters.band[23] ;
 wire \filters.band[24] ;
 wire \filters.band[25] ;
 wire \filters.band[26] ;
 wire \filters.band[27] ;
 wire \filters.band[28] ;
 wire \filters.band[29] ;
 wire \filters.band[2] ;
 wire \filters.band[30] ;
 wire \filters.band[31] ;
 wire \filters.band[3] ;
 wire \filters.band[4] ;
 wire \filters.band[5] ;
 wire \filters.band[6] ;
 wire \filters.band[7] ;
 wire \filters.band[8] ;
 wire \filters.band[9] ;
 wire \filters.bp ;
 wire \filters.cutoff_lut[10] ;
 wire \filters.cutoff_lut[11] ;
 wire \filters.cutoff_lut[12] ;
 wire \filters.cutoff_lut[13] ;
 wire \filters.cutoff_lut[14] ;
 wire \filters.cutoff_lut[15] ;
 wire \filters.cutoff_lut[16] ;
 wire \filters.cutoff_lut[6] ;
 wire \filters.cutoff_lut[7] ;
 wire \filters.cutoff_lut[8] ;
 wire \filters.cutoff_lut[9] ;
 wire \filters.filt_1 ;
 wire \filters.filt_2 ;
 wire \filters.filt_3 ;
 wire \filters.filter_step[0] ;
 wire \filters.filter_step[1] ;
 wire \filters.filter_step[2] ;
 wire \filters.high[0] ;
 wire \filters.high[10] ;
 wire \filters.high[11] ;
 wire \filters.high[12] ;
 wire \filters.high[13] ;
 wire \filters.high[14] ;
 wire \filters.high[15] ;
 wire \filters.high[16] ;
 wire \filters.high[17] ;
 wire \filters.high[18] ;
 wire \filters.high[19] ;
 wire \filters.high[1] ;
 wire \filters.high[20] ;
 wire \filters.high[21] ;
 wire \filters.high[22] ;
 wire \filters.high[23] ;
 wire \filters.high[24] ;
 wire \filters.high[25] ;
 wire \filters.high[26] ;
 wire \filters.high[27] ;
 wire \filters.high[28] ;
 wire \filters.high[29] ;
 wire \filters.high[2] ;
 wire \filters.high[30] ;
 wire \filters.high[31] ;
 wire \filters.high[3] ;
 wire \filters.high[4] ;
 wire \filters.high[5] ;
 wire \filters.high[6] ;
 wire \filters.high[7] ;
 wire \filters.high[8] ;
 wire \filters.high[9] ;
 wire \filters.hp ;
 wire \filters.low[0] ;
 wire \filters.low[10] ;
 wire \filters.low[11] ;
 wire \filters.low[12] ;
 wire \filters.low[13] ;
 wire \filters.low[14] ;
 wire \filters.low[15] ;
 wire \filters.low[16] ;
 wire \filters.low[17] ;
 wire \filters.low[18] ;
 wire \filters.low[19] ;
 wire \filters.low[1] ;
 wire \filters.low[20] ;
 wire \filters.low[21] ;
 wire \filters.low[22] ;
 wire \filters.low[23] ;
 wire \filters.low[24] ;
 wire \filters.low[25] ;
 wire \filters.low[26] ;
 wire \filters.low[27] ;
 wire \filters.low[28] ;
 wire \filters.low[29] ;
 wire \filters.low[2] ;
 wire \filters.low[30] ;
 wire \filters.low[31] ;
 wire \filters.low[3] ;
 wire \filters.low[4] ;
 wire \filters.low[5] ;
 wire \filters.low[6] ;
 wire \filters.low[7] ;
 wire \filters.low[8] ;
 wire \filters.low[9] ;
 wire \filters.lp ;
 wire \filters.mode_vol[0] ;
 wire \filters.mode_vol[1] ;
 wire \filters.mode_vol[2] ;
 wire \filters.mode_vol[3] ;
 wire \filters.mode_vol[7] ;
 wire \filters.res_filt[3] ;
 wire \filters.res_filt[4] ;
 wire \filters.res_filt[5] ;
 wire \filters.res_filt[6] ;
 wire \filters.res_filt[7] ;
 wire \filters.res_lut[0] ;
 wire \filters.res_lut[10] ;
 wire \filters.res_lut[1] ;
 wire \filters.res_lut[2] ;
 wire \filters.res_lut[3] ;
 wire \filters.res_lut[4] ;
 wire \filters.res_lut[5] ;
 wire \filters.res_lut[6] ;
 wire \filters.res_lut[7] ;
 wire \filters.res_lut[8] ;
 wire \filters.res_lut[9] ;
 wire \filters.sample_buff[0] ;
 wire \filters.sample_buff[10] ;
 wire \filters.sample_buff[11] ;
 wire \filters.sample_buff[12] ;
 wire \filters.sample_buff[13] ;
 wire \filters.sample_buff[14] ;
 wire \filters.sample_buff[1] ;
 wire \filters.sample_buff[2] ;
 wire \filters.sample_buff[3] ;
 wire \filters.sample_buff[4] ;
 wire \filters.sample_buff[5] ;
 wire \filters.sample_buff[6] ;
 wire \filters.sample_buff[7] ;
 wire \filters.sample_buff[8] ;
 wire \filters.sample_buff[9] ;
 wire \filters.sample_filtered[0] ;
 wire \filters.sample_filtered[10] ;
 wire \filters.sample_filtered[11] ;
 wire \filters.sample_filtered[12] ;
 wire \filters.sample_filtered[13] ;
 wire \filters.sample_filtered[14] ;
 wire \filters.sample_filtered[15] ;
 wire \filters.sample_filtered[1] ;
 wire \filters.sample_filtered[2] ;
 wire \filters.sample_filtered[3] ;
 wire \filters.sample_filtered[4] ;
 wire \filters.sample_filtered[5] ;
 wire \filters.sample_filtered[6] ;
 wire \filters.sample_filtered[7] ;
 wire \filters.sample_filtered[8] ;
 wire \filters.sample_filtered[9] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net8;
 wire net9;
 wire \spi_dac_i.counter[0] ;
 wire \spi_dac_i.counter[1] ;
 wire \spi_dac_i.counter[2] ;
 wire \spi_dac_i.counter[3] ;
 wire \spi_dac_i.counter[4] ;
 wire \spi_dac_i.spi_dat_buff_0[0] ;
 wire \spi_dac_i.spi_dat_buff_0[10] ;
 wire \spi_dac_i.spi_dat_buff_0[11] ;
 wire \spi_dac_i.spi_dat_buff_0[1] ;
 wire \spi_dac_i.spi_dat_buff_0[2] ;
 wire \spi_dac_i.spi_dat_buff_0[3] ;
 wire \spi_dac_i.spi_dat_buff_0[4] ;
 wire \spi_dac_i.spi_dat_buff_0[5] ;
 wire \spi_dac_i.spi_dat_buff_0[6] ;
 wire \spi_dac_i.spi_dat_buff_0[7] ;
 wire \spi_dac_i.spi_dat_buff_0[8] ;
 wire \spi_dac_i.spi_dat_buff_0[9] ;
 wire \spi_dac_i.spi_dat_buff_1[0] ;
 wire \spi_dac_i.spi_dat_buff_1[10] ;
 wire \spi_dac_i.spi_dat_buff_1[11] ;
 wire \spi_dac_i.spi_dat_buff_1[1] ;
 wire \spi_dac_i.spi_dat_buff_1[2] ;
 wire \spi_dac_i.spi_dat_buff_1[3] ;
 wire \spi_dac_i.spi_dat_buff_1[4] ;
 wire \spi_dac_i.spi_dat_buff_1[5] ;
 wire \spi_dac_i.spi_dat_buff_1[6] ;
 wire \spi_dac_i.spi_dat_buff_1[7] ;
 wire \spi_dac_i.spi_dat_buff_1[8] ;
 wire \spi_dac_i.spi_dat_buff_1[9] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[0].attenuation.in ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[1].attenuation.in ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[2].attenuation.in ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ;
 wire \tt_um_rejunity_sn76489.chan[3].attenuation.in ;
 wire \tt_um_rejunity_sn76489.clk_counter[0] ;
 wire \tt_um_rejunity_sn76489.clk_counter[1] ;
 wire \tt_um_rejunity_sn76489.clk_counter[2] ;
 wire \tt_um_rejunity_sn76489.clk_counter[3] ;
 wire \tt_um_rejunity_sn76489.clk_counter[4] ;
 wire \tt_um_rejunity_sn76489.control_noise[0][0] ;
 wire \tt_um_rejunity_sn76489.control_noise[0][1] ;
 wire \tt_um_rejunity_sn76489.control_noise[0][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][0] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][1] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][3] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][4] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][5] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][6] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][7] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][8] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[0][9] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][0] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][1] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][3] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][4] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][5] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][6] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][7] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][8] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[1][9] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][0] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][1] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][2] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][3] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][4] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][5] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][6] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][7] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][8] ;
 wire \tt_um_rejunity_sn76489.control_tone_freq[2][9] ;
 wire \tt_um_rejunity_sn76489.latch_control_reg[0] ;
 wire \tt_um_rejunity_sn76489.latch_control_reg[1] ;
 wire \tt_um_rejunity_sn76489.latch_control_reg[2] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.restart_noise ;
 wire \tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[7] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[8] ;
 wire \tt_um_rejunity_sn76489.tone[0].gen.counter[9] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[7] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[8] ;
 wire \tt_um_rejunity_sn76489.tone[1].gen.counter[9] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[0] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[1] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[2] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[3] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[4] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[5] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[6] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[7] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[8] ;
 wire \tt_um_rejunity_sn76489.tone[2].gen.counter[9] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A2 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A1 (.I(\filters.res_filt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A1 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A2 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A1 (.I(\filters.res_filt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A1 (.I(\filters.res_filt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A1 (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A1 (.I(\filters.res_filt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A1 (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A1 (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__A1 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__I (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__A1 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__I (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__I (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A1 (.I(\clk_trg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__A1 (.I(\clk_trg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__I (.I(\clk_trg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__I (.I(\clk_trg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__A1 (.I(\channels.clk_div[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__A2 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__A1 (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__A2 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__S1 (.I(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__I (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__I (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__A1 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__B1 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__B2 (.I(\channels.ring_outs[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__I (.I(\channels.clk_div[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__A2 (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__I (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__A1 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__A2 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__I (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__A2 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__B1 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__B2 (.I(\channels.ring_outs[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__I (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__I (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__I (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__I (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__I (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__I (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__I (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08675__I (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__I (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__I (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__I (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__I (.I(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__I (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__I (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__I (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__I (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__I (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__I (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__I (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__I (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__I (.I(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__I (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__I (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__S0 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__S1 (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__I (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__I (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__I (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__I (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__S1 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__A2 (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__S1 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__S1 (.I(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__A1 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__S0 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__S1 (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__I (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__I (.I(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A2 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A2 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A2 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__A2 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__B2 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__I (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A2 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A2 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A2 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__I (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__I (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A1 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A2 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__I (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__B1 (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__B2 (.I(\channels.ring_outs[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__I (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A2 (.I(\channels.ctrl_reg2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A2 (.I(\channels.ctrl_reg3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__B1 (.I(\channels.ctrl_reg1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A1 (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A1 (.I(\channels.ctrl_reg3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A2 (.I(\channels.sync_outs[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A3 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A1 (.I(\channels.ctrl_reg2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A2 (.I(\channels.sync_outs[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A3 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A1 (.I(\channels.ctrl_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A2 (.I(\channels.sync_outs[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__I (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A1 (.I(\channels.freq3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A1 (.I(\channels.freq2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__B2 (.I(\channels.freq1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__I (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__I (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__I (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__A1 (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A1 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A1 (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__C (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A1 (.I(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A1 (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__I (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__I (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A1 (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A2 (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__I (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__I (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A1 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__C (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A1 (.I(\channels.freq3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A1 (.I(\channels.freq2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__B2 (.I(\channels.freq1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__I (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__S0 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__S1 (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A1 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__A2 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A1 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A1 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__A1 (.I(\channels.freq3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__A1 (.I(\channels.freq2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__B2 (.I(\channels.freq1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__S0 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__S1 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A1 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A1 (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A1 (.I(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A1 (.I(\channels.freq3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__A1 (.I(\channels.freq2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__B2 (.I(\channels.freq1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__S0 (.I(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__S1 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A1 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__I (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A1 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A1 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__S0 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__S1 (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A1 (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A1 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A1 (.I(\channels.freq3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__B2 (.I(\channels.freq1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__S0 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__S1 (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A1 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A1 (.I(\channels.freq2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__B2 (.I(\channels.freq1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__S0 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__S1 (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A1 (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A1 (.I(\channels.freq3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A1 (.I(\channels.freq2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__B2 (.I(\channels.freq1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__S0 (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__S1 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A1 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__A2 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__A1 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__I (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A1 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A1 (.I(\channels.freq2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__B2 (.I(\channels.freq1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__S0 (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__S1 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A1 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__A1 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__A2 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A1 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A2 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__A1 (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__I (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__B1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__I (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A1 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__A1 (.I(\channels.freq2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__B2 (.I(\channels.freq1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__S0 (.I(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__S1 (.I(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__I (.I(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A1 (.I(\channels.freq3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A1 (.I(\channels.freq2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__B2 (.I(\channels.freq1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__S1 (.I(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A1 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__B1 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A1 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A1 (.I(\channels.freq3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A1 (.I(\channels.freq2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__B2 (.I(\channels.freq1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__I (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A2 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__A1 (.I(\channels.freq2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__B2 (.I(\channels.freq1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__S0 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__S1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__I (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A2 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__B1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A2 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__A1 (.I(\channels.freq2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__B2 (.I(\channels.freq1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__I (.I(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__S1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__I (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A2 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A2 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A1 (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A2 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A1 (.I(\channels.freq2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__B2 (.I(\channels.freq1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__S0 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__S1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__I (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A1 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__B1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A2 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A1 (.I(\channels.freq3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A1 (.I(\channels.freq2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__B2 (.I(\channels.freq1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A1 (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A2 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__I (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A2 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A2 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__I (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A1 (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A2 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__B (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__S0 (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__S1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__I (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09076__A3 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__B (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__I (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__B1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__S0 (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__S1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__I (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__A1 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__A2 (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A1 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__A2 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__S0 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__S1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__I (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A1 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A2 (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__B (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A1 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A2 (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A3 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A1 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__B1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__I (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__S0 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__S1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__I (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__I (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A2 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A2 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A1 (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__B1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A3 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__S0 (.I(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__S1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__I (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A2 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A2 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A1 (.I(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__I (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A2 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__S0 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__S1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A2 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__A1 (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__B1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A2 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A1 (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A2 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__S0 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__S1 (.I(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__S0 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__S1 (.I(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A1 (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A2 (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__I (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__A1 (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__A3 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__I (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__I (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A1 (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A2 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__S0 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__S1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__B1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__I (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__I (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__I (.I(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__I (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__I (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__S0 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__S1 (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__B1 (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__I (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__S0 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__S1 (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__B1 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__I (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__I (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__I (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__S0 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__S1 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__S0 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__S1 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__I (.I(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__S0 (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__S1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__B1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__I (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__S0 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__S1 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__S0 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__S1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__B1 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__S0 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__S1 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__B2 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__I (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__I (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__S0 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__S1 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__B2 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__I (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__I (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__S0 (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__S1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__B1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__B2 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__S0 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__S1 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__B2 (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__S0 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__S1 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__B2 (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__I3 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__S0 (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__S1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__B1 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__B2 (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__S0 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__S1 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__B1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__B2 (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__S0 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__S1 (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__B1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__B2 (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__S1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A1 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__I (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A1 (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A2 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A1 (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__I (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__I (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__I (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A1 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__I (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__I (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__I (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__I (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A1 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__I (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__I (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A1 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09344__A1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__I (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__I (.I(\filters.filt_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__I (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__I (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__B (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A1 (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09367__I (.I(\filters.filt_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__I (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__I (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__I (.I(\filters.filt_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__A1 (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__I (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A1 (.I(\filters.res_filt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__I (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__I (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__I (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__A2 (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A1 (.I(\filters.mode_vol[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A1 (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A1 (.I(\filters.mode_vol[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A1 (.I(\filters.mode_vol[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__I (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A1 (.I(\filters.lp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A1 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__I (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__I (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__A1 (.I(\filters.bp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__B (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__I (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__I (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__A1 (.I(\filters.hp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__B (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__I (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__I (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__A1 (.I(\filters.mode_vol[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__B (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__I (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__I (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A1 (.I(\channels.ctrl_reg2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A2 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A1 (.I(\channels.atk_dec2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A2 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__B1 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__B2 (.I(\channels.pw3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__I (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__I (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__A1 (.I(\filters.cutoff_lut[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__B1 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A1 (.I(\channels.freq1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__B2 (.I(\channels.ctrl_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__A1 (.I(\channels.sus_rel3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__B1 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__B2 (.I(\channels.pw2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A2 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__B2 (.I(\channels.pw2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__I (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__I (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A1 (.I(\channels.atk_dec3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A2 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__B2 (.I(\channels.sus_rel2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__C1 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__C2 (.I(\channels.freq3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A3 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__I (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__I (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A1 (.I(\channels.ch3_env[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__I (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A1 (.I(\channels.freq2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A2 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__B2 (.I(\channels.ctrl_reg3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__I (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__A1 (.I(\channels.pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__B2 (.I(\channels.freq1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A1 (.I(\channels.pw1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__B2 (.I(\channels.freq2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__A1 (.I(\filters.mode_vol[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__B2 (.I(\channels.pw3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A2 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__A1 (.I(\channels.sample3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__B2 (.I(\clk_trg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__I (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__B1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A1 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A1 (.I(\channels.ctrl_reg2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A2 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A1 (.I(\channels.atk_dec2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A2 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__B1 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__B2 (.I(\channels.pw3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A1 (.I(\filters.cutoff_lut[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__B1 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__B2 (.I(\filters.cutoff_lut[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A1 (.I(\channels.freq1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__B2 (.I(\channels.ctrl_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A1 (.I(\channels.sus_rel3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__B2 (.I(\channels.pw2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A1 (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A2 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__B2 (.I(\channels.pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(\channels.atk_dec3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A2 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__B2 (.I(\channels.sus_rel2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__C1 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__C2 (.I(\channels.freq3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__A3 (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A1 (.I(\channels.ch3_env[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A1 (.I(\channels.freq2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A2 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__B2 (.I(\channels.ctrl_reg3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A1 (.I(\channels.pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__B2 (.I(\channels.freq1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__A1 (.I(\channels.pw1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__B2 (.I(\channels.freq2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A1 (.I(\filters.mode_vol[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A2 (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__B2 (.I(\channels.pw3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A2 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A1 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__B2 (.I(\clk_trg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__B1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A1 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__I (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__I (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__I (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A1 (.I(\channels.ctrl_reg3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__B1 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__B2 (.I(\channels.pw2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__I (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__I (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A1 (.I(\channels.sus_rel2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__B2 (.I(\channels.freq3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A1 (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A2 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A1 (.I(\channels.pw1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__B1 (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__B2 (.I(\channels.ctrl_reg1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A1 (.I(\filters.cutoff_lut[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__B2 (.I(\channels.sus_rel3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__A1 (.I(\channels.sus_rel1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__A2 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__B2 (.I(\channels.sample3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A1 (.I(\channels.atk_dec1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A1 (.I(\channels.pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A2 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__B2 (.I(\channels.freq2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__A1 (.I(\channels.ctrl_reg2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__B2 (.I(\channels.freq2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A1 (.I(\channels.pw3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__B2 (.I(\channels.pw2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A1 (.I(\channels.ch3_env[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A2 (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__B2 (.I(\channels.freq1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A1 (.I(\filters.cutoff_lut[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A2 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__B2 (.I(\channels.atk_dec3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__A1 (.I(\channels.atk_dec2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__B2 (.I(\channels.pw3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A1 (.I(\channels.freq1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A2 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__B2 (.I(\channels.freq3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A1 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A1 (.I(\channels.sus_rel3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__B1 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__B2 (.I(\channels.sus_rel1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(\filters.res_filt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A2 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__B2 (.I(\channels.freq2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A1 (.I(\filters.mode_vol[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A2 (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__B1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__B2 (.I(\channels.sus_rel2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A1 (.I(\channels.ch3_env[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__B2 (.I(\channels.pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__A1 (.I(\channels.pw3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__B1 (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__B2 (.I(\channels.freq1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A1 (.I(\channels.atk_dec2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(\channels.pw1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A1 (.I(\channels.freq3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__B2 (.I(\channels.freq2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A1 (.I(\channels.ctrl_reg1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A2 (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__B2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A1 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__A1 (.I(\channels.ctrl_reg2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__B2 (.I(\channels.ctrl_reg3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A1 (.I(\channels.pw2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A2 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__B2 (.I(\channels.atk_dec1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A1 (.I(\channels.atk_dec3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A2 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__B2 (.I(\channels.pw3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A1 (.I(\filters.cutoff_lut[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A2 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__B2 (.I(\channels.freq1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A1 (.I(\channels.freq3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__B1 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__B2 (.I(\channels.pw2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A1 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__I (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A1 (.I(\filters.cutoff_lut[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A1 (.I(\channels.sus_rel3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__B2 (.I(\channels.freq1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__I (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A1 (.I(\channels.ctrl_reg2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__B2 (.I(\channels.atk_dec2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__I (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A1 (.I(\channels.pw2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__B2 (.I(\channels.freq2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__I (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__B2 (.I(\channels.ctrl_reg3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__I (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__I (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__B2 (.I(\channels.ctrl_reg1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__I (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A1 (.I(\filters.res_filt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__B2 (.I(\channels.sample3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A1 (.I(\channels.ch3_env[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__B2 (.I(\channels.atk_dec1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A1 (.I(\filters.lp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__B1 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__B2 (.I(\channels.sus_rel1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A2 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__B (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A2 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__A1 (.I(\filters.cutoff_lut[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A1 (.I(\channels.sus_rel3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__B1 (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__B2 (.I(\channels.freq1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A1 (.I(\channels.ctrl_reg2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A1 (.I(\channels.pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__B2 (.I(\channels.freq2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A1 (.I(\channels.freq3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A2 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__A1 (.I(\channels.pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__B2 (.I(\channels.ctrl_reg1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__A1 (.I(\filters.res_filt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__B2 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A1 (.I(\channels.ch3_env[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__B2 (.I(\channels.atk_dec1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__A1 (.I(\channels.freq1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__B2 (.I(\channels.pw3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A1 (.I(\filters.bp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__B1 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__B2 (.I(\channels.sus_rel1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__I (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A2 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__B (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A2 (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__A1 (.I(\filters.cutoff_lut[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A1 (.I(\channels.sus_rel3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__B1 (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__B2 (.I(\channels.freq1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A1 (.I(\channels.ctrl_reg2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__A1 (.I(\channels.pw2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__B2 (.I(\channels.freq2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__A2 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__B1 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__B2 (.I(\channels.freq2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A1 (.I(\channels.pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__B2 (.I(\channels.ctrl_reg1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A1 (.I(\filters.res_filt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__B2 (.I(\channels.sample3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__A1 (.I(\channels.ch3_env[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__B2 (.I(\channels.atk_dec1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A1 (.I(\channels.freq1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__B2 (.I(\channels.pw3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__A1 (.I(\filters.hp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__B1 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__B2 (.I(\channels.sus_rel1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__B (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__A2 (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A1 (.I(\filters.mode_vol[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A2 (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__B2 (.I(\channels.freq3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__I (.I(\channels.sample3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A1 (.I(\channels.ctrl_reg2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A2 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__B2 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__A1 (.I(\channels.atk_dec1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A4 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__A1 (.I(\channels.ch3_env[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__B1 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__B2 (.I(\channels.sus_rel1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A1 (.I(\channels.freq1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A2 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A1 (.I(\channels.atk_dec3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__B2 (.I(\channels.freq2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A1 (.I(\channels.freq2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__B2 (.I(\channels.freq1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A1 (.I(\channels.atk_dec2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A2 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__B2 (.I(\channels.freq3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__B2 (.I(\channels.ctrl_reg1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__A1 (.I(\filters.cutoff_lut[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__B2 (.I(\channels.sus_rel3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A1 (.I(\filters.res_filt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__B2 (.I(\channels.pw3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(\channels.pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__B2 (.I(\channels.pw2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__B (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A2 (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A1 (.I(\channels.freq1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__B (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A1 (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A1 (.I(\channels.freq1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A1 (.I(\channels.freq1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(\channels.freq1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A1 (.I(\channels.freq1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A1 (.I(\channels.freq1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__A1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A1 (.I(\channels.freq1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__A1 (.I(\channels.freq1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__I (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__A1 (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A1 (.I(\channels.pw1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__A1 (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A1 (.I(\channels.pw1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__B (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A1 (.I(\channels.pw1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__B (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A1 (.I(\channels.pw1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__B (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__I (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A2 (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__I (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__I (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A1 (.I(\channels.ctrl_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__B (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__I (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__I (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__A1 (.I(\channels.ctrl_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__A1 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__I (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__A1 (.I(\channels.ctrl_reg1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A1 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__I (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__A1 (.I(\channels.ctrl_reg1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__I (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__I (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__A1 (.I(\channels.ctrl_reg1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__A1 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__A1 (.I(\channels.ctrl_reg1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__A1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A1 (.I(\channels.ctrl_reg1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A1 (.I(\channels.ctrl_reg1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A1 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__A1 (.I(\channels.atk_dec1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A1 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A1 (.I(\channels.atk_dec1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__A1 (.I(\channels.atk_dec1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A1 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__A1 (.I(\channels.atk_dec1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__A1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__A1 (.I(\channels.atk_dec1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A1 (.I(\channels.atk_dec1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__I (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__I (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__A1 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A1 (.I(\channels.sus_rel1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__A1 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A1 (.I(\channels.sus_rel1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__I (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A1 (.I(\channels.sus_rel1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__I (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A1 (.I(\channels.sus_rel1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__I (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(\channels.sus_rel1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__I (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A1 (.I(\channels.sus_rel1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A1 (.I(\channels.freq2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__A1 (.I(\channels.freq2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A1 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A1 (.I(\channels.freq2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__A1 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A1 (.I(\channels.freq2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__A1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__A1 (.I(\channels.freq2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A1 (.I(\channels.freq2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__B (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A1 (.I(\channels.freq2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__B (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__A1 (.I(\channels.freq2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__B (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__I (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A1 (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A2 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__I (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__I (.I(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A1 (.I(\channels.pw2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__B (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__I (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__I (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A1 (.I(\channels.pw2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__A1 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__I (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__I (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__A1 (.I(\channels.pw2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__I (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A1 (.I(\channels.pw2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__A2 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__A1 (.I(\channels.ctrl_reg2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__A1 (.I(\channels.ctrl_reg2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__A1 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A1 (.I(\channels.ctrl_reg2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__A1 (.I(\channels.ctrl_reg2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A1 (.I(\channels.ctrl_reg2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__A1 (.I(\channels.ctrl_reg2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__A1 (.I(\channels.ctrl_reg2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A1 (.I(\channels.ctrl_reg2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__A2 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A1 (.I(\channels.atk_dec2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__A1 (.I(\channels.atk_dec2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A1 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A1 (.I(\channels.atk_dec2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A1 (.I(\channels.atk_dec2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A1 (.I(\channels.atk_dec2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__I (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__I (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__A1 (.I(\channels.atk_dec2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__I (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__I (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__I (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A1 (.I(\channels.sus_rel2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__I (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__A1 (.I(\channels.sus_rel2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__B (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__A1 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__A1 (.I(\channels.sus_rel2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__B (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A1 (.I(\channels.sus_rel2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__B (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__I (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__I (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__B (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__A1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__I (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__I (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__I (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__I (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A1 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__I (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A2 (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__A1 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__I (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__I (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A1 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__I (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A1 (.I(\channels.freq3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A1 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__I (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__A1 (.I(\channels.freq3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__A1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__I (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A1 (.I(\channels.freq3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A1 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A1 (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__A1 (.I(\channels.pw3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__A1 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A1 (.I(\channels.pw3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__A1 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A1 (.I(\channels.pw3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A1 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A1 (.I(\channels.pw3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__A2 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__A1 (.I(\channels.ctrl_reg3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A1 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A1 (.I(\channels.ctrl_reg3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__A1 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A1 (.I(\channels.ctrl_reg3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__A1 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A1 (.I(\channels.ctrl_reg3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A1 (.I(\channels.ctrl_reg3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__B (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__B (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__B (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A1 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__A2 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__A1 (.I(\channels.atk_dec3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__B (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__A1 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__I (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__I (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__A1 (.I(\channels.atk_dec3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__A1 (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__A1 (.I(\channels.atk_dec3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A1 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__A1 (.I(\channels.atk_dec3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__I (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__B (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__B (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__A1 (.I(\channels.atk_dec3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__B (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__A1 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__I (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__I (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__I (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__I (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__A1 (.I(\channels.sus_rel3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__B (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__I (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__I (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__A1 (.I(\channels.sus_rel3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A1 (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__I (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__A1 (.I(\channels.sus_rel3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A1 (.I(\channels.sus_rel3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__I (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__I (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A1 (.I(\channels.sus_rel3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A1 (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__I (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__I (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__A1 (.I(\channels.sus_rel3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__A1 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__I (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__A1 (.I(\channels.sus_rel3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__I (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A1 (.I(\channels.sus_rel3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__A1 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A2 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__I (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__I (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__I (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__I (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A1 (.I(\filters.cutoff_lut[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__A1 (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A1 (.I(\filters.cutoff_lut[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__A1 (.I(\filters.cutoff_lut[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__I (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__I (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__A1 (.I(\filters.cutoff_lut[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__A1 (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__I (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__A1 (.I(\filters.cutoff_lut[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__A1 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A1 (.I(\filters.cutoff_lut[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A1 (.I(\filters.cutoff_lut[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__A1 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__I (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A1 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__I (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__A2 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__I (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__A2 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__C (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A2 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__A2 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__C (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A1 (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A2 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__I (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__I (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A1 (.I(\channels.sync_outs[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A1 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__I (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__A1 (.I(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__A2 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__I (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__A1 (.I(\channels.sync_outs[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__A2 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A1 (.I(\channels.sync_outs[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A2 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__A2 (.I(\channels.ctrl_reg2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A2 (.I(\channels.ctrl_reg3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__B1 (.I(\channels.ctrl_reg1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A1 (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__I (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A1 (.I(\channels.ctrl_reg2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A2 (.I(\channels.ring_outs[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A1 (.I(\channels.ctrl_reg3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A2 (.I(\channels.ring_outs[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A1 (.I(\channels.ctrl_reg1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A2 (.I(\channels.ring_outs[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__I (.I(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A1 (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__A1 (.I(\channels.ctrl_reg1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__B2 (.I(\channels.ctrl_reg2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__I (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__A1 (.I(\channels.ctrl_reg2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__B2 (.I(\channels.ctrl_reg1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__I (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A1 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__A1 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__A3 (.I(\channels.pw3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A2 (.I(\channels.pw2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__A1 (.I(\channels.pw1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__A3 (.I(\channels.pw2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__A3 (.I(\channels.pw3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A1 (.I(\channels.pw1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__S0 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__S1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__A1 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__B2 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__I (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__A2 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__A3 (.I(\channels.pw3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__A2 (.I(\channels.pw2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__A1 (.I(\channels.pw1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A3 (.I(\channels.pw2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A2 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A3 (.I(\channels.pw3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A1 (.I(\channels.pw1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__B2 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__A1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A1 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__B2 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__B2 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__A3 (.I(\channels.pw2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__A3 (.I(\channels.pw3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__A1 (.I(\channels.pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A1 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__I (.I(\channels.pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A2 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A3 (.I(\channels.pw3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__A2 (.I(\channels.pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__C (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A2 (.I(\channels.pw2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__C (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__A3 (.I(\channels.pw2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A2 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A3 (.I(\channels.pw3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A1 (.I(\channels.pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A3 (.I(\channels.pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__A1 (.I(\channels.pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__A1 (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A1 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__C2 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__I (.I(\channels.pw2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__A2 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__A3 (.I(\channels.pw3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__A1 (.I(\channels.pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A3 (.I(\channels.pw2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A2 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A3 (.I(\channels.pw3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A1 (.I(\channels.pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A1 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A3 (.I(\channels.pw3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__A2 (.I(\channels.pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__A2 (.I(\channels.pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__A1 (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__B (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__I (.I(\channels.pw2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A2 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A3 (.I(\channels.pw3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__A1 (.I(\channels.pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__A1 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__B2 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A3 (.I(\channels.pw2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__A1 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__A1 (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__B (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__A2 (.I(\channels.ctrl_reg2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__B1 (.I(\channels.ctrl_reg1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A1 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__I (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__I2 (.I(\channels.ch3_env[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__S0 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__S1 (.I(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__I (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A1 (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A2 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A1 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__I (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A1 (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A2 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__I (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__I (.I(\channels.ch3_env[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__I (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A3 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__I (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__I (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__I (.I(\channels.ch3_env[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A1 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__I (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__I2 (.I(\channels.ch3_env[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__A2 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__A3 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A2 (.I(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__I (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A1 (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A2 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__A1 (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A1 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__I (.I(\channels.ch3_env[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A1 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A1 (.I(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__S (.I(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A1 (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A1 (.I(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__I (.I(\channels.ch3_env[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A2 (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__S (.I(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__I (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A2 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__I (.I(\channels.ch3_env[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A2 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A2 (.I(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A2 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A2 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A1 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__I (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__I (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__A2 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__I (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__I (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__A3 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__I (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__A1 (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__A2 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__A2 (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__A1 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__I (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__I (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__I (.I(\channels.ch3_env[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__A1 (.I(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__A2 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A2 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A3 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__I (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__A1 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__A2 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A2 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A3 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__A2 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__I (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A2 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__A3 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A1 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__A3 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__A2 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__A1 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__I (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A3 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__A3 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__A3 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__I (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__A1 (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A1 (.I(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__A2 (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__A3 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__I (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__I (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__A2 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__B1 (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A2 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__A1 (.I(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A1 (.I(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__A2 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A2 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__A1 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__A3 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A2 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A3 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A1 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__A2 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__A1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A1 (.I(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A3 (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__A1 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__A1 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__A1 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__A2 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A1 (.I(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__A1 (.I(\channels.sample3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A1 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A2 (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__A1 (.I(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__A1 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A2 (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__A1 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__A1 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__A2 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__A1 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__I (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__A1 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__A2 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10575__A1 (.I(\channels.sample3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__A1 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__A2 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__I (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__I (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__A1 (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__A3 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__B1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__A4 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__A2 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10605__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__A1 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__A1 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__I (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A1 (.I(\channels.sample3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__A1 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__A2 (.I(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__A2 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A1 (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A3 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__A2 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A1 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__A1 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__A1 (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__A1 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A1 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__A1 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__A2 (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__A1 (.I(\channels.sample3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__I (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__A1 (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A1 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A2 (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__A1 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__A2 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__A1 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__I (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__A2 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A1 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A2 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__I (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__A1 (.I(\channels.sample3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__A2 (.I(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A1 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__I (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__A1 (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__A1 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__A2 (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A1 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__A1 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__A1 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__I (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__A2 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A2 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__I (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A1 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__A1 (.I(\channels.sample3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A2 (.I(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A2 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__A1 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10831__A2 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A2 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__A2 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__I (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__A1 (.I(\channels.sample3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__A2 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__A2 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__A1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__A2 (.I(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A1 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A2 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__A1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A1 (.I(\channels.sample3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__A2 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A1 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__A1 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__A2 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__I (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A1 (.I(\channels.sample2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A2 (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A1 (.I(\channels.sample2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A1 (.I(\channels.sample2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A2 (.I(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A1 (.I(\channels.sample2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__I (.I(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__A1 (.I(\channels.sample2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A2 (.I(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A1 (.I(\channels.sample2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(\channels.sample2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A2 (.I(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A1 (.I(\channels.sample2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__A2 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__I (.I(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A1 (.I(\channels.sample2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A2 (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A2 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A1 (.I(\channels.sample2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A2 (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A2 (.I(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A1 (.I(\channels.sample2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A2 (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A2 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A1 (.I(\channels.sample2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A2 (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A1 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A2 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__I (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A1 (.I(\channels.sample1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A2 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A2 (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__I (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A1 (.I(\channels.sample1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__A1 (.I(\channels.sample1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A2 (.I(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A1 (.I(\channels.sample1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__A1 (.I(\channels.sample1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A2 (.I(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__I (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A1 (.I(\channels.sample1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A2 (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A1 (.I(\channels.sample1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A2 (.I(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A1 (.I(\channels.sample1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__A2 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A1 (.I(\channels.sample1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A2 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A1 (.I(\channels.sample1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__A2 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__A2 (.I(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A1 (.I(\channels.sample1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A2 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__A2 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A1 (.I(\channels.sample1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A2 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__A2 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__I (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__I (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__I (.I(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__I (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__A1 (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__A1 (.I(\filters.low[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__B (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__A2 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__A1 (.I(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__I (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__I (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__I (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__I (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A1 (.I(\filters.lp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A2 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A1 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A1 (.I(\filters.hp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A2 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__B2 (.I(\filters.bp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__C (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A3 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__B1 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__B (.I(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__A2 (.I(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__B (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A1 (.I(\filters.high[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__A1 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__B1 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__B2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__B (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__I (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__B (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__A1 (.I(\filters.high[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__B (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__B (.I(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__A1 (.I(\filters.high[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__B (.I(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__A1 (.I(\filters.low[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__B (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__I (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__B (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A1 (.I(\filters.high[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__B (.I(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__I (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A1 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__B (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A1 (.I(\filters.high[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__I (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A2 (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__B (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__B (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__I (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__A1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__B (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__A2 (.I(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__I (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__I (.I(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__B (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__A1 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__A2 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__B (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__A1 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A2 (.I(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__I (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__B (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__A1 (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__B (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__A1 (.I(\filters.high[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__B (.I(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__B (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A1 (.I(\filters.high[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__A1 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__A1 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__B1 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__A1 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A1 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A2 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A1 (.I(\filters.high[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__A1 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A2 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A1 (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__I (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__I (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__I (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__I (.I(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__B (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__A2 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A1 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__B1 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A1 (.I(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A2 (.I(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A1 (.I(\filters.cutoff_lut[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__I (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__A1 (.I(\filters.cutoff_lut[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11283__A1 (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__A1 (.I(\filters.cutoff_lut[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11291__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__I (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__A2 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A1 (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A2 (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__I (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__I (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__A1 (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__I (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__I (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__I (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__C (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A1 (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__I (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__I (.I(\tt_um_rejunity_sn76489.control_tone_freq[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__A1 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__I (.I(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__I (.I(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__A1 (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__C (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__I (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__A1 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__I (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__A1 (.I(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__I (.I(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__I (.I(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__I (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__B (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A1 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__B (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A1 (.I(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__B (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__A1 (.I(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__S0 (.I(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__S1 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11346__I (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__S0 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__S1 (.I(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__I (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__I (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A1 (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A2 (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__A1 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__I (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__A1 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11360__A1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A3 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11363__A1 (.I(\channels.ctrl_reg2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11363__A2 (.I(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11364__A1 (.I(\channels.ctrl_reg3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11364__A2 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11364__B2 (.I(\channels.ctrl_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__A1 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11368__I (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__A1 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__B (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__A3 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__A4 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__I (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__A2 (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__A1 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__A2 (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A1 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A2 (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__A1 (.I(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__I (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__A2 (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__A1 (.I(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__I (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__B1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__I (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__A1 (.I(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__B1 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__A1 (.I(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__B1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__A1 (.I(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__B1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__I (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11416__I (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__I (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__B1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A2 (.I(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__B1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__B1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__B1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__I (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__I (.I(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11438__A2 (.I(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11439__A1 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A2 (.I(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__A1 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__A2 (.I(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11447__A1 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__I (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__A2 (.I(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A1 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__I (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__I (.I(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__B1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__I (.I(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__A1 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__B1 (.I(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__A1 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__B1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11467__A1 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__B1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__I (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__I (.I(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11475__I (.I(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11476__B1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__A2 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__B2 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11480__B1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__B1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__B1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__A2 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__A1 (.I(\channels.freq1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__B (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11498__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11500__A1 (.I(\channels.freq1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__A1 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11502__A1 (.I(\channels.freq1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__A1 (.I(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11504__A1 (.I(\channels.freq1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__A1 (.I(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11510__I (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__A2 (.I(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__I (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__I (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__I (.I(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__B (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__A1 (.I(\channels.freq1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__A1 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__A2 (.I(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__A1 (.I(\channels.freq1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11521__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11521__A2 (.I(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__A1 (.I(\channels.freq1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__A1 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__A2 (.I(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__I (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__A2 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11530__A1 (.I(\channels.pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11531__A1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11533__A1 (.I(\channels.pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11534__A1 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A1 (.I(\channels.pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11537__A1 (.I(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__A1 (.I(\channels.pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11539__A1 (.I(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__A1 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11542__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11543__C (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11544__A1 (.I(\channels.pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__A1 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__A1 (.I(\channels.pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11547__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11549__I (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__A1 (.I(\channels.pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__A1 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11553__A2 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__A1 (.I(\channels.freq2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__A1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__A1 (.I(\channels.freq2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__A1 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__I (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11563__A1 (.I(\channels.freq2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__A1 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11566__A1 (.I(\channels.freq2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11567__A1 (.I(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__B (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__I (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11575__A1 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__I (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__A1 (.I(\channels.freq2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__I (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__A1 (.I(\channels.freq2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11581__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11587__A1 (.I(\channels.freq3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11588__A1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__A1 (.I(\channels.freq3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11590__A1 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11591__A1 (.I(\channels.freq3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11592__A1 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11594__A1 (.I(\channels.freq3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11600__B (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A1 (.I(\channels.freq3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11603__A1 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__A1 (.I(\channels.freq3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11607__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__A1 (.I(\channels.pw3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11613__A1 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11614__I (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__A1 (.I(\channels.pw3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11617__A1 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__A1 (.I(\channels.pw3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11619__A1 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11620__A1 (.I(\channels.pw3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__B (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11627__A1 (.I(\channels.pw3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11628__A1 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__A1 (.I(\channels.pw3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11631__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__A1 (.I(\channels.pw3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11633__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11635__A2 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11639__A1 (.I(\channels.pw2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__A1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11641__A1 (.I(\channels.pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__A1 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__A1 (.I(\channels.pw2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11645__A1 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__A1 (.I(\channels.pw2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11647__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11649__A1 (.I(\channels.pw2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11649__A2 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11650__I (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11652__A1 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__I (.I(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__B (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11655__A1 (.I(\channels.pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11656__A1 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11657__A1 (.I(\channels.pw2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11658__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__A1 (.I(\channels.pw2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__B (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11661__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__A2 (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11665__I (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11666__I (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11667__I (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__I (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11669__I (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__A1 (.I(\channels.clk_div[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__B (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11671__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__I (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11673__A1 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11673__A2 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11674__I (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__A1 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11677__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__A1 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11681__I (.I(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__I (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11684__I (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11685__I (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11686__I (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11687__I (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11691__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11693__A1 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11695__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11696__I (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11697__A1 (.I(\channels.sus_rel1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__A1 (.I(\channels.sus_rel3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__A2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__A2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__A1 (.I(\channels.sus_rel1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11702__A1 (.I(\channels.sus_rel3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__I0 (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__S (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11704__A1 (.I(\channels.sus_rel3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__B2 (.I(\channels.sus_rel1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11706__A1 (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11707__A1 (.I(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11708__A1 (.I(\channels.sus_rel3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11709__B2 (.I(\channels.sus_rel1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__B1 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__A2 (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__B1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__B2 (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11713__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11713__B1 (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11713__B2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__A2 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__A1 (.I(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__A2 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11717__A2 (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11717__B1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11717__B2 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__A1 (.I(\channels.sus_rel3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__B2 (.I(\channels.sus_rel2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11723__I (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11724__I (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11725__A1 (.I(\channels.atk_dec3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11725__B2 (.I(\channels.atk_dec2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11726__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11728__S (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11730__I (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11731__B2 (.I(\channels.atk_dec2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11731__C2 (.I(\channels.atk_dec1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11734__A1 (.I(\channels.atk_dec3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11734__B2 (.I(\channels.atk_dec2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11735__A1 (.I(\channels.sus_rel3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11735__B2 (.I(\channels.sus_rel2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11737__S (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11738__A2 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11738__B (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11739__C2 (.I(\channels.atk_dec1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11741__I (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11743__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11744__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11745__A1 (.I(\channels.sus_rel3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11745__B2 (.I(\channels.sus_rel2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11746__A1 (.I(\channels.atk_dec3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11746__B2 (.I(\channels.atk_dec2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11747__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11748__I0 (.I(\channels.atk_dec1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11748__I1 (.I(\channels.sus_rel1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11748__S (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11750__C2 (.I(\channels.atk_dec1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11753__I (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__A1 (.I(\channels.atk_dec3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__B2 (.I(\channels.atk_dec2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11757__A1 (.I(\channels.sus_rel3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11757__B2 (.I(\channels.sus_rel2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11758__S (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11759__I0 (.I(\channels.atk_dec1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11759__I1 (.I(\channels.sus_rel1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11761__A1 (.I(\channels.atk_dec3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11761__B2 (.I(\channels.atk_dec2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11761__C2 (.I(\channels.atk_dec1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11763__I (.I(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11765__A1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11765__A2 (.I(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11767__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__I (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11771__I (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__S0 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__S1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11774__I (.I(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11776__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11777__A2 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11781__I (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11782__S0 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11782__S1 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__I (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11789__I (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11793__S0 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11793__S1 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11800__S0 (.I(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11800__S1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__S0 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__S1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11807__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__S0 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__S1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11814__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11818__S0 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11818__S1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11822__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11826__S0 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11826__S1 (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11831__S0 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11831__S1 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__S0 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__S0 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__S1 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11843__A2 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11844__S0 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11844__S1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11847__A1 (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__S0 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__S1 (.I(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11853__I (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11855__S (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11857__A1 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11858__A1 (.I(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11858__C (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11859__A1 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11864__S0 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11864__S1 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11865__A2 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11866__A2 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11868__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11869__A2 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11874__I (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11875__A2 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11876__I (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11877__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__I (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11879__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11879__B (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11884__A2 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11885__I (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11891__I (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11902__I (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11909__A2 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11911__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11922__A1 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__A2 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11932__A1 (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11941__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11949__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11949__A2 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11950__A1 (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11952__A1 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__I (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11955__I (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11957__A1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11958__I (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11962__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11967__I (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11969__A1 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11977__I (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11979__A1 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11980__I (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11989__A1 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11992__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11993__B (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11994__A1 (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11996__A2 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11997__I (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11998__I (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12001__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__I (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12006__A1 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12012__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12018__A1 (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12022__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12027__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12031__A1 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12031__B (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12032__A1 (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12035__A1 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12036__I (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12038__A1 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__I (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12041__A2 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12043__A2 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__A2 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__A2 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12049__I (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12050__I (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12058__A1 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12059__I (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12060__I (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__A2 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__A3 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12080__I (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12082__A1 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12082__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12083__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12084__I (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12086__A1 (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12087__I (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12097__I (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12098__I (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12106__A1 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12107__I (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12108__I (.I(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__A1 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__B (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12128__A1 (.I(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12128__B (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12181__I (.I(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12182__A1 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12182__A2 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12183__I (.I(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__A4 (.I(\filters.high[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12187__I (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12188__A1 (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12188__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12194__A2 (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12195__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12197__I (.I(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12200__A4 (.I(\filters.high[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12201__A1 (.I(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12201__A2 (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__A1 (.I(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12207__A1 (.I(\filters.res_lut[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12208__I (.I(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__I (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12210__I (.I(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12213__I (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12215__A1 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12215__A2 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12215__A3 (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12216__A4 (.I(\filters.high[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12220__A1 (.I(\filters.res_lut[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12221__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12222__I (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12223__I (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12224__A1 (.I(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12224__A3 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12229__A1 (.I(\filters.res_lut[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12230__I (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12233__I (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12239__A1 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12239__A3 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12240__I (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12241__I (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12242__I0 (.I(\filters.cutoff_lut[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12243__I (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12244__I (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12245__I (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12247__I (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12248__A1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12248__A3 (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12249__A4 (.I(\filters.high[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12250__I (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12253__I (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12255__I (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12257__A3 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12259__I (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12260__I (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12262__A3 (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12263__I0 (.I(\filters.cutoff_lut[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12267__A1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12267__A3 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12268__A4 (.I(\filters.high[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12272__A1 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12272__A3 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12281__I (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12283__I (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12284__A3 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12286__A1 (.I(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12288__A1 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12291__I (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12292__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12292__A2 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12295__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12296__A1 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12296__A3 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12297__A1 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12297__A2 (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12301__I (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12303__A2 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12305__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12306__I (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12309__A1 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12309__A2 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12314__I (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12318__I (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12319__I (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12320__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12321__I (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12323__B2 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12324__A1 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12324__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12324__A3 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12326__I (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12335__A1 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12339__I (.I(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12340__I (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12341__I (.I(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12343__A1 (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12343__A2 (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12344__A2 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12347__I0 (.I(\filters.cutoff_lut[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12348__I (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12349__I (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12351__A1 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12352__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12352__A2 (.I(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12356__I (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12360__I (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12361__A2 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12365__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12366__A4 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12367__I (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12368__I (.I(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12369__A1 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12369__A2 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12369__A3 (.I(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12370__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12370__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12370__A3 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12379__I (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12380__I (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12382__A2 (.I(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12385__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12391__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12391__A2 (.I(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12392__I (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12394__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12396__A1 (.I(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12397__A1 (.I(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12398__I0 (.I(\filters.cutoff_lut[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12399__I (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12400__I (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12401__I (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12405__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12409__I (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12411__A2 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12415__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12416__I (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12418__A1 (.I(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12420__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12423__A1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12423__A2 (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12424__A1 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12425__A4 (.I(\filters.high[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12427__A1 (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12427__A2 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12429__I (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12430__A1 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12430__A2 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12465__A1 (.I(\filters.cutoff_lut[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12467__I (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12471__A1 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12471__A2 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12472__I (.I(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12473__I (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12474__I (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12475__I (.I(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12476__I (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12477__A1 (.I(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12477__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12477__B1 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12478__A2 (.I(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12480__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12481__A3 (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12482__A1 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12482__A2 (.I(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12484__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12485__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12489__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12489__A2 (.I(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12489__A3 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12490__I (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12491__I (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12493__A2 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12494__A3 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12495__A2 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12496__I (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12498__A1 (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12499__I (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12501__I (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12503__A1 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12505__A2 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12507__A1 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12508__I (.I(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12509__A4 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12510__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12511__I (.I(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12513__A1 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12515__A1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12515__A2 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12520__A2 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12522__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12525__I (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12526__I (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12528__A1 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12528__B1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12529__A4 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12533__I (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12534__A1 (.I(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12543__I (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12544__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12545__A1 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12547__A1 (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12547__A2 (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12547__A3 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12551__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12551__A2 (.I(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12556__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12561__A1 (.I(\filters.res_lut[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12562__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12569__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12582__I (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12583__A1 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12583__A2 (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12585__I (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12586__A1 (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12586__A2 (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12586__A3 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12588__A2 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12588__A3 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12592__I (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12593__A1 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12593__A2 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12596__A1 (.I(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12597__I (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12600__A2 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12601__I (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__A3 (.I(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12604__A1 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12606__A2 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12608__A1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12609__A1 (.I(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12611__A1 (.I(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12612__A1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12615__A2 (.I(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12618__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12618__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12619__I (.I(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12620__I (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12621__A1 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12621__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12622__I (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12623__I (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12624__I (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12625__A1 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12625__B2 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12626__A1 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12626__A2 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12626__A4 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12628__A1 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12628__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12632__A1 (.I(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12634__A1 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12636__A1 (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12636__A2 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12637__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12639__I (.I(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12641__I (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12642__A2 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12642__A3 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12642__A4 (.I(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12643__I (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12644__A2 (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12646__A1 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12654__I (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12656__I (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12657__I (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12658__A1 (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12658__A2 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12658__A4 (.I(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12659__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12660__I (.I(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12661__A1 (.I(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12661__A2 (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12662__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12662__B2 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12663__A2 (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12664__I (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12665__A2 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12666__I (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12667__I (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12668__I (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12670__I (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12671__A2 (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12673__A1 (.I(\filters.res_lut[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12673__A2 (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12674__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12674__B2 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12675__A2 (.I(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12678__A1 (.I(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12681__I0 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12690__A1 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12691__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12692__I (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12693__A1 (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12703__A1 (.I(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12703__A2 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12707__A2 (.I(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12707__A3 (.I(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12707__B (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12721__I (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12722__B2 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12723__I (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12724__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12724__A2 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12727__I (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12729__I (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12730__A1 (.I(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12732__A1 (.I(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12732__A2 (.I(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12733__A1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12734__I (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12735__I0 (.I(\filters.high[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12735__S (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12736__I (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12737__I (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12738__A1 (.I(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12740__A2 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12742__A1 (.I(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12742__A2 (.I(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12745__A3 (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12746__I (.I(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12747__I (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12748__A1 (.I(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12748__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12749__A1 (.I(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12749__A2 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12749__A3 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12756__A1 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12756__A2 (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12757__A1 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12757__A3 (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12761__A1 (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12763__I (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12764__A1 (.I(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12764__A2 (.I(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12765__S (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12766__I (.I(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12767__A1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12767__A2 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12768__A2 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12770__A1 (.I(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12770__A2 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12775__I (.I(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12776__I (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12777__I (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12779__A1 (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12779__A2 (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12784__I (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12785__A1 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12788__I (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12791__I (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12792__I (.I(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12794__I (.I(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12795__A1 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12796__A1 (.I(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12798__A2 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12799__A2 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12805__A1 (.I(\filters.cutoff_lut[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12805__A2 (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12807__A1 (.I(\filters.cutoff_lut[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12809__I (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12810__A1 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12810__A3 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12811__A1 (.I(\filters.cutoff_lut[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12812__I (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12813__A3 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12814__A1 (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12815__A1 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12816__A1 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12816__A2 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12817__A1 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12817__A2 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12818__A1 (.I(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12820__I (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12821__A3 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12822__A2 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12823__A3 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12824__A2 (.I(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12824__A3 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12826__A1 (.I(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12826__A2 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12828__A2 (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12829__I (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12830__I (.I(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12833__A1 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12833__B2 (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12834__A1 (.I(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12834__A2 (.I(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12841__A1 (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12842__A1 (.I(\filters.cutoff_lut[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12843__I (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12845__I (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12847__A1 (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12847__A2 (.I(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12848__A3 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12849__A3 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12850__I (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12852__A3 (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12854__A1 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12854__A2 (.I(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12858__A1 (.I(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12859__A1 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12860__A1 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12861__A1 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12864__A1 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12864__A2 (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12864__A3 (.I(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12867__A1 (.I(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12867__A2 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12869__A1 (.I(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12869__A2 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12871__A1 (.I(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12871__A2 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12873__I (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12875__A1 (.I(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12875__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12875__B2 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12877__A1 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12877__A2 (.I(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12879__A1 (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12880__I (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12881__A2 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12882__A3 (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12883__A1 (.I(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12884__I (.I(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12885__A2 (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12886__I0 (.I(\filters.high[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12886__S (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12887__I (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12889__A1 (.I(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12889__A2 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12890__A1 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12890__A2 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12891__A2 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12892__A1 (.I(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12903__A1 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12903__A2 (.I(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12904__A1 (.I(\filters.cutoff_lut[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12908__A1 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12908__A2 (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12909__I (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12910__A2 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12910__A3 (.I(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12912__A3 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12913__A3 (.I(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12916__A1 (.I(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12916__A2 (.I(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12918__A4 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12921__A1 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12921__A2 (.I(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12925__A1 (.I(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12926__A2 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12927__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12927__A2 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12927__A3 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12928__A1 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12928__A2 (.I(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12930__A1 (.I(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12930__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12930__A3 (.I(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12932__A1 (.I(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12934__A1 (.I(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12936__A1 (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12936__A2 (.I(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12937__A1 (.I(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12937__A2 (.I(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12938__A1 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12941__A1 (.I(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12942__A1 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12942__A2 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12943__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12944__A1 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12947__I (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12948__A2 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12949__S (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12950__I (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12951__A1 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12951__A2 (.I(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12952__A2 (.I(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12958__A1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12959__A1 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12964__A1 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12965__A1 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12967__I (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12969__A2 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12972__A2 (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12975__A1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12975__A2 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12977__A1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12977__A2 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12979__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12980__A1 (.I(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12980__A2 (.I(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12984__A2 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12987__A1 (.I(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12991__A1 (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12992__A1 (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12997__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13015__A1 (.I(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13015__A2 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13020__A1 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13022__A2 (.I(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13024__A2 (.I(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13047__A3 (.I(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13057__A1 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13058__A2 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13064__A1 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13076__A2 (.I(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13077__I (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13078__A1 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13078__A2 (.I(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13080__A1 (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13084__A1 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13084__A2 (.I(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13085__A1 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13085__A2 (.I(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13086__A1 (.I(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13087__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13087__B1 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13087__B2 (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13088__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13088__A2 (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13088__A4 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13090__A1 (.I(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13090__A2 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13091__A1 (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13091__A2 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13091__A3 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13093__A2 (.I(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13093__A3 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13094__A2 (.I(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13096__A1 (.I(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13097__I (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13099__A2 (.I(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13100__I1 (.I(\filters.band[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13101__I (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13103__A1 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13103__A2 (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13104__A1 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13104__A2 (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13110__A2 (.I(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13116__A1 (.I(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13116__A2 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13125__A1 (.I(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13125__A2 (.I(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13127__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13127__A3 (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13128__A2 (.I(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13129__A1 (.I(\filters.cutoff_lut[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13131__A1 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13131__A2 (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13133__A2 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13135__A3 (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13138__A2 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13139__A1 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13139__A2 (.I(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13141__A2 (.I(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13146__A1 (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13147__A2 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13148__A3 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13149__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13151__A2 (.I(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13157__A2 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13163__A2 (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13172__A2 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13173__A2 (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13176__A1 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13176__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13177__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13181__A2 (.I(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13182__A1 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13183__A1 (.I(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13183__A3 (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13184__A2 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13187__A2 (.I(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13188__A1 (.I(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13190__A1 (.I(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13192__A1 (.I(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13193__A1 (.I(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13195__A2 (.I(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13197__A2 (.I(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13198__A1 (.I(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13203__A1 (.I(\filters.band[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13204__A2 (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13205__A2 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13206__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13207__I (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13208__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13209__S (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13210__I (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13212__A1 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13212__A2 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13213__A1 (.I(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13213__A2 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13223__A1 (.I(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13225__A2 (.I(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13226__A1 (.I(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13228__A1 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13228__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13229__I (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13230__A1 (.I(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13230__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13235__A1 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13237__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13240__A1 (.I(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13240__A2 (.I(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13241__A2 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13251__I (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13253__A2 (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13254__A3 (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13257__A1 (.I(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13258__A3 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13259__A2 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13259__A3 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13260__A2 (.I(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13262__A2 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13267__A1 (.I(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13268__A1 (.I(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13270__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13270__B2 (.I(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13271__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13271__A2 (.I(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13271__A4 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13273__A2 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13274__A1 (.I(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13274__A2 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13275__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13275__A2 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13278__A2 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13279__A1 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13279__A2 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13280__I1 (.I(\filters.band[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13280__S (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13281__I (.I(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13282__A1 (.I(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13283__A1 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13284__A2 (.I(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13289__I (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13290__A2 (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13291__A2 (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13296__A1 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13296__A2 (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13297__A1 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13298__A1 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13299__A1 (.I(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13303__A2 (.I(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13325__A1 (.I(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13325__A2 (.I(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13329__A1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13329__A2 (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13330__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13335__A2 (.I(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__A3 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__A4 (.I(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13337__A2 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13337__B1 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13338__A3 (.I(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13339__A2 (.I(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13341__A2 (.I(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13344__A2 (.I(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13345__I (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13346__A1 (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13346__A3 (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13348__A1 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13348__A2 (.I(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13349__A2 (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13350__A1 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13358__A1 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13359__A1 (.I(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13361__B1 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13362__A1 (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13362__A2 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13362__A4 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13364__A2 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13365__A2 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13366__A1 (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13366__A2 (.I(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13368__A1 (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13368__A2 (.I(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13369__I (.I(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13370__A1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13370__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13371__A1 (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13371__A2 (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13372__S (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13373__I (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13374__A1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13376__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13377__A1 (.I(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13381__A1 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13381__A2 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13387__A1 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13387__A2 (.I(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13388__A1 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13389__I (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13392__A1 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13392__A3 (.I(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13395__A1 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13397__A2 (.I(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13399__A2 (.I(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13402__A1 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13402__A2 (.I(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13407__A1 (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13428__A1 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13428__A2 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13432__A1 (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13440__A1 (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13440__A2 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13445__A1 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13445__A2 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13447__A3 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13448__A1 (.I(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13448__A2 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13449__A1 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13449__A2 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13451__A1 (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13451__A2 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13452__A1 (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13452__A2 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13452__B1 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13452__B2 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13454__A1 (.I(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13454__A2 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13456__A1 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13456__A2 (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13460__A2 (.I(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13462__A2 (.I(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13464__A1 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13464__A2 (.I(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13464__A3 (.I(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13468__A1 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13469__I (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13471__A1 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13471__A3 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13473__A1 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13476__A1 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13486__I (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13489__A1 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13489__A3 (.I(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13490__A2 (.I(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13491__I (.I(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13492__A1 (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13492__A2 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13493__A1 (.I(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13494__I (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13495__A1 (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13500__A1 (.I(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13500__B (.I(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13501__A1 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13502__A1 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13502__A2 (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13502__A3 (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13503__A1 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13508__A2 (.I(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13514__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13514__A2 (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13519__I (.I(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13520__A2 (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13521__A2 (.I(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13526__A1 (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13527__A2 (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13528__I1 (.I(\filters.band[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13529__I (.I(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13530__A1 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13531__A1 (.I(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13535__I (.I(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13536__A1 (.I(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13536__B1 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13536__B2 (.I(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13537__A1 (.I(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13537__A2 (.I(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13537__A4 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13539__A1 (.I(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13541__A1 (.I(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13541__A2 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13543__A1 (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13544__A1 (.I(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13545__A1 (.I(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13549__A3 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13553__A1 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13553__A2 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13555__I (.I(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13556__I (.I(\filters.low[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13557__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13557__A2 (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13562__I (.I(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13563__B (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13564__A1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13565__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13566__I (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13568__I (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13569__I (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13571__A1 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13571__A2 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13573__A2 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13574__A2 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13576__A1 (.I(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13582__I (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13584__A1 (.I(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13585__I (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13586__A1 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13588__A1 (.I(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13593__A2 (.I(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13594__A1 (.I(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13595__A1 (.I(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13595__A2 (.I(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13602__I (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13604__A1 (.I(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13607__A1 (.I(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13608__A1 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13609__I1 (.I(\filters.band[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13610__A2 (.I(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13613__I (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13614__A1 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13614__B1 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13614__B2 (.I(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13615__A1 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13615__A2 (.I(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13617__A1 (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13617__A2 (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13619__A1 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13619__A2 (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13620__A2 (.I(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13620__A3 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13621__A1 (.I(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13623__A1 (.I(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13633__A1 (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13634__A1 (.I(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13634__A2 (.I(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13635__A1 (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13639__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13639__A2 (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13641__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13642__A1 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13642__A3 (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13643__A1 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13643__A2 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13648__I (.I(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13649__A2 (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13649__B1 (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13651__I (.I(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13655__A2 (.I(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13656__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13656__A2 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13658__A2 (.I(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13658__A3 (.I(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13659__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13668__A1 (.I(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13669__A3 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13670__B (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13673__A1 (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13674__A1 (.I(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13674__A2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13677__A1 (.I(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13678__A1 (.I(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13678__C (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13679__A1 (.I(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13679__A2 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13680__A1 (.I(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13681__A1 (.I(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13683__C (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13688__I (.I(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13689__A1 (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13690__A1 (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13692__A1 (.I(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13695__A1 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13698__A1 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13698__A2 (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13700__A1 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13700__A2 (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13708__A1 (.I(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13711__A1 (.I(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13711__A2 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13714__I (.I(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13715__A1 (.I(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13716__A1 (.I(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13717__I1 (.I(\filters.band[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13718__A2 (.I(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13721__A1 (.I(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13721__A2 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13722__A1 (.I(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13722__A2 (.I(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13725__A2 (.I(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13726__A1 (.I(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13728__A3 (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13729__A1 (.I(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13739__A1 (.I(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13740__A2 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13741__A1 (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13742__A2 (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13745__A1 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13747__A2 (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13749__A1 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13749__A2 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13750__A1 (.I(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13750__A2 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13751__A2 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13753__A1 (.I(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13753__A2 (.I(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13754__A1 (.I(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13754__A2 (.I(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13756__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13757__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13758__A1 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13758__A2 (.I(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13761__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13761__A2 (.I(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13765__A2 (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13772__A1 (.I(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13772__A2 (.I(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13773__A1 (.I(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13774__A2 (.I(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13776__I (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13778__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13779__A2 (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13785__A1 (.I(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13786__C (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13792__I (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13793__A1 (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13794__A1 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13796__A1 (.I(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13802__A2 (.I(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13804__A1 (.I(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13804__A2 (.I(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13809__A1 (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13810__A1 (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13812__I (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13816__A1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13816__A2 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13819__I (.I(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13820__A1 (.I(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13821__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13822__I1 (.I(\filters.band[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13823__A2 (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13826__A1 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13826__A2 (.I(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13826__B1 (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13826__B2 (.I(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13827__A1 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13827__A2 (.I(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13827__A3 (.I(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13827__A4 (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13828__A2 (.I(_05828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13829__A1 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13830__A1 (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13830__A2 (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13831__A1 (.I(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13833__A1 (.I(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13833__A2 (.I(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13835__A1 (.I(_05820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13839__A1 (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13840__A1 (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13842__A2 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13843__A2 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13845__A2 (.I(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13846__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13847__A1 (.I(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13851__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13851__A2 (.I(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13853__A2 (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13856__A1 (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13856__A2 (.I(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13860__A1 (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13861__A3 (.I(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13862__A1 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13862__A3 (.I(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13869__A2 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13869__A3 (.I(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13874__A1 (.I(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13874__A2 (.I(_05875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13875__A1 (.I(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13875__A2 (.I(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13877__A1 (.I(_05878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13877__A2 (.I(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13878__I (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13879__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13880__A1 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13881__A1 (.I(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13888__A1 (.I(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13889__A1 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13889__C (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13890__A1 (.I(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13891__A1 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13892__A1 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13894__A2 (.I(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13896__A2 (.I(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13897__A3 (.I(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13898__A2 (.I(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13898__A3 (.I(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13899__A1 (.I(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13899__A2 (.I(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13900__A1 (.I(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13900__A2 (.I(_05875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13901__A1 (.I(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13901__A2 (.I(_05875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13909__I (.I(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13910__A1 (.I(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13910__A2 (.I(_05910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13911__A1 (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13913__A1 (.I(_05820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13916__A1 (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13916__A2 (.I(_05910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13918__A1 (.I(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13921__A1 (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13926__A1 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13926__A2 (.I(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13927__A1 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13927__A2 (.I(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13929__A1 (.I(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13929__A2 (.I(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13931__A1 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13931__A2 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13934__A1 (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13934__A2 (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13935__A1 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13935__A2 (.I(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13936__I1 (.I(\filters.band[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13936__S (.I(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13937__A1 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13937__A2 (.I(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13942__A4 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13944__A1 (.I(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13947__A1 (.I(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13949__A1 (.I(_05944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13949__A2 (.I(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13951__A1 (.I(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13959__B2 (.I(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13960__A2 (.I(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13962__A1 (.I(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13964__A2 (.I(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13972__A2 (.I(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13973__A2 (.I(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13974__A1 (.I(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13974__A2 (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13979__A1 (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13984__A2 (.I(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13984__A3 (.I(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13992__A1 (.I(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13992__A2 (.I(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13993__I (.I(\filters.low[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13994__A1 (.I(_05994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13995__A1 (.I(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13996__A1 (.I(_05993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13998__B (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13999__A1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14000__I (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14007__A1 (.I(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14007__A2 (.I(_06006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14008__I (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14009__A1 (.I(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14009__A2 (.I(_05910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14011__A1 (.I(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14015__I (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14019__A1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14024__A1 (.I(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14024__A2 (.I(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14025__A1 (.I(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14025__A2 (.I(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14027__A1 (.I(_05944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14027__A2 (.I(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14031__I (.I(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14032__A1 (.I(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14033__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14033__A2 (.I(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14034__I0 (.I(\filters.high[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14034__S (.I(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14035__A1 (.I(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14035__A2 (.I(_06034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14038__A1 (.I(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14039__A1 (.I(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14039__A3 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14041__A1 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14041__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14042__A1 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14043__A2 (.I(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14044__A1 (.I(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14045__A1 (.I(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14047__A1 (.I(_06030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14053__A1 (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14054__A2 (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14056__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14057__A2 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14059__A1 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14059__A2 (.I(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14061__A1 (.I(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14062__A1 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14062__A2 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14063__A1 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14063__A2 (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14067__A2 (.I(_06066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14071__A1 (.I(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14071__A2 (.I(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14072__A3 (.I(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14074__A1 (.I(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14075__A1 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14078__A1 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14081__A1 (.I(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14081__A2 (.I(_06080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14089__A1 (.I(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14089__A2 (.I(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14089__B (.I(_06088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14090__A1 (.I(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14093__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14093__A2 (.I(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14094__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14094__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14095__A1 (.I(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14096__A1 (.I(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14098__I (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14099__A1 (.I(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14099__A2 (.I(_06098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14099__B (.I(_05993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14105__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14106__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14114__A1 (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14115__A1 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14115__A2 (.I(_06006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14118__A1 (.I(_06030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14119__A1 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14121__A1 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14123__A1 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14128__A1 (.I(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14128__A2 (.I(_06080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14130__A2 (.I(_06066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14132__A1 (.I(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14137__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14139__A1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14142__A1 (.I(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14142__A2 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14143__A1 (.I(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14145__A2 (.I(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14155__A1 (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14155__A2 (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14156__A1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14156__A2 (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14157__A1 (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14157__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14162__A1 (.I(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14162__A2 (.I(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14163__A1 (.I(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14168__A1 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14169__A1 (.I(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14169__A2 (.I(_06034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14170__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14170__A2 (.I(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14171__A1 (.I(\filters.band[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14171__A2 (.I(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14174__A1 (.I(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14175__A1 (.I(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14177__A1 (.I(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14177__A2 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14178__A1 (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14178__A2 (.I(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14180__A2 (.I(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14184__A1 (.I(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14195__A1 (.I(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14195__A2 (.I(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14199__A1 (.I(_06088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14200__I (.I(_06198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14201__A1 (.I(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14202__A1 (.I(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14204__A1 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14205__A1 (.I(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14205__A2 (.I(_06202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14206__A2 (.I(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14212__A1 (.I(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14218__A1 (.I(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14218__A2 (.I(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14230__A1 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14231__A1 (.I(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14231__A2 (.I(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14233__A2 (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14236__A1 (.I(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14238__A1 (.I(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14238__A2 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14239__A1 (.I(_06234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14239__A2 (.I(_06235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14248__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14249__A1 (.I(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14255__A1 (.I(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14255__A2 (.I(_06252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14262__A1 (.I(\filters.band[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14262__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14263__A1 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14264__A1 (.I(\filters.band[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14264__A2 (.I(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14268__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14269__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14271__A1 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14275__A1 (.I(_06259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14279__I (.I(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14282__A1 (.I(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14284__A1 (.I(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14287__I (.I(_06034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14288__A1 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14290__A1 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14292__A1 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14304__A1 (.I(_06299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14304__A2 (.I(_06301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14305__I (.I(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14308__B (.I(_06305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14310__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14311__A2 (.I(_06202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14312__A2 (.I(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14314__A2 (.I(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14315__A2 (.I(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14322__A2 (.I(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14323__A2 (.I(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14323__B2 (.I(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14326__A1 (.I(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14328__A1 (.I(_06299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14328__A2 (.I(_06301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14329__A1 (.I(_06305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14329__B2 (.I(_06198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14330__A1 (.I(_06299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14330__A2 (.I(_06301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14331__A1 (.I(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14336__A1 (.I(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14336__A2 (.I(_06252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14347__A1 (.I(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14347__A2 (.I(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14348__A1 (.I(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14354__A1 (.I(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14355__A1 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14357__A2 (.I(_06353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14359__A1 (.I(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14359__A2 (.I(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14361__A1 (.I(_06234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14361__A2 (.I(_06235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14362__A1 (.I(_06234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14362__A2 (.I(_06235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14366__A1 (.I(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14373__A1 (.I(_06338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14373__A2 (.I(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14380__A1 (.I(\filters.band[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14380__A2 (.I(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14381__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14388__I (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14389__A1 (.I(_06385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14390__A1 (.I(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14395__A1 (.I(_06376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14400__A1 (.I(_06259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14406__I (.I(\filters.band[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14407__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14410__A1 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14410__A2 (.I(_06406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14416__A1 (.I(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14421__A2 (.I(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14424__A1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14424__A2 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14425__A1 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14425__A2 (.I(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14426__A1 (.I(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14426__A2 (.I(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14429__A1 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14430__I (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14437__A1 (.I(_06338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14437__A2 (.I(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14444__A2 (.I(_06353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14448__A2 (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14449__A1 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14449__A2 (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14450__A1 (.I(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14452__A1 (.I(_06443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14456__A1 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14459__A2 (.I(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14461__I (.I(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14462__A1 (.I(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14462__A2 (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14467__A1 (.I(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14468__A1 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14469__A1 (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14472__A1 (.I(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14482__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14483__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14483__A2 (.I(_06034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14484__A2 (.I(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14489__A1 (.I(_06385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14490__A1 (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14490__A2 (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14501__A1 (.I(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14502__A1 (.I(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14502__A2 (.I(_06406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14504__A1 (.I(_06376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14507__A2 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14511__I (.I(\filters.band[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14512__A2 (.I(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14519__A1 (.I(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14522__A2 (.I(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14527__A1 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14527__A2 (.I(_06202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14528__A1 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14528__A2 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14529__A1 (.I(_06522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14529__A2 (.I(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14530__A1 (.I(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14530__A2 (.I(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14535__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14536__A1 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14550__A1 (.I(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14556__A2 (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14560__A2 (.I(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14571__A1 (.I(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14574__A1 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14574__A2 (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14576__A1 (.I(\filters.band[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14581__A1 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14584__A1 (.I(_06385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14585__A1 (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14591__A2 (.I(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14594__A1 (.I(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14594__A2 (.I(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14596__A1 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14599__A1 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14600__A1 (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14605__A1 (.I(_06443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14609__A1 (.I(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14614__A1 (.I(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14615__A1 (.I(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14615__A2 (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14616__A1 (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14616__A2 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14617__A2 (.I(_06610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14621__A2 (.I(_06615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14622__A2 (.I(_06615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14631__A2 (.I(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14632__A1 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14632__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14633__A1 (.I(_06625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14633__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14635__A1 (.I(_06522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14635__A2 (.I(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14636__A1 (.I(_06522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14636__A2 (.I(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14641__A1 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14646__A1 (.I(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14647__A1 (.I(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14649__A1 (.I(_06385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14653__A1 (.I(\filters.band[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14655__A1 (.I(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14655__A2 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14656__A1 (.I(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14656__A2 (.I(_06406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14660__A1 (.I(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14664__A1 (.I(_06610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14665__A1 (.I(_06610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14667__A1 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14668__A1 (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14668__A2 (.I(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14673__A1 (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14673__A2 (.I(_06006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14676__A1 (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14676__A2 (.I(_06406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14678__A3 (.I(_06671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14682__A1 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14682__A2 (.I(_05910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14683__A1 (.I(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14683__A2 (.I(_06006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14685__A1 (.I(\filters.band[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14686__A1 (.I(_06676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14686__A2 (.I(_06678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14687__A1 (.I(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14694__A1 (.I(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14695__A1 (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14695__A2 (.I(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14696__A1 (.I(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14700__A1 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14701__A2 (.I(_06693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14712__A2 (.I(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14719__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14719__A2 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14720__A1 (.I(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14720__A2 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14721__A1 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14721__A2 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14722__A1 (.I(_06625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14722__A2 (.I(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14725__B (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14726__A1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14732__A1 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14732__A2 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14734__A2 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14737__A1 (.I(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14737__A2 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14740__I (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14741__A2 (.I(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14742__A2 (.I(_06733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14743__A1 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14745__I (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14746__I (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14747__B (.I(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14748__A1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14751__I (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14754__A1 (.I(_06745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14756__A1 (.I(_06747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14758__A2 (.I(_06733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14759__A1 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14759__A2 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14760__A1 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14763__A1 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14764__A1 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14764__A2 (.I(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14765__A1 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14765__A2 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14769__B (.I(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14773__A1 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14775__A2 (.I(_06733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14776__A2 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14778__A1 (.I(_06747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14783__I (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14784__C (.I(_06773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14785__I (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14788__B (.I(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14792__I (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14793__I0 (.I(\filters.low[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14793__I1 (.I(\filters.band[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14793__S (.I(_06781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14796__A1 (.I(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14797__I (.I(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14798__I (.I(_06786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14799__A1 (.I(\filters.band[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14799__B (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14802__I (.I(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14806__A1 (.I(_06793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14808__I0 (.I(\filters.low[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14808__S (.I(_06781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14811__B (.I(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14813__I (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14814__I1 (.I(\filters.band[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14814__S (.I(_06098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14816__B (.I(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14820__A1 (.I(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14821__I (.I(_06786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14822__A1 (.I(\filters.band[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14822__A2 (.I(_06808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14822__B (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14824__S (.I(_06781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14825__A1 (.I(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14827__A1 (.I(_06793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14829__A1 (.I(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14830__A2 (.I(_06808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14830__B (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14832__I1 (.I(\filters.band[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14832__S (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14833__A1 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14836__B (.I(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14840__A1 (.I(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14841__I (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14843__A1 (.I(\filters.band[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14843__A2 (.I(_06808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14845__I (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14847__A1 (.I(_06793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14848__I1 (.I(\filters.band[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14848__S (.I(_06098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14849__A1 (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14852__A1 (.I(\filters.band[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14852__A2 (.I(_06808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14854__I0 (.I(\filters.low[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14854__I1 (.I(\filters.band[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14854__S (.I(_06098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14857__B (.I(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14861__I (.I(_06786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14862__A1 (.I(\filters.band[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14865__A1 (.I(\filters.band[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14865__A2 (.I(_06781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14866__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14868__A1 (.I(_06745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14872__A1 (.I(\filters.band[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14876__B (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14879__I (.I(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14881__A1 (.I(\filters.band[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14883__A1 (.I(_06860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14885__A1 (.I(\filters.band[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14885__B (.I(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14888__A1 (.I(_06747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14889__A1 (.I(_06859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14890__S (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14891__A1 (.I(_06860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14897__I (.I(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14898__I (.I(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14899__I1 (.I(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14899__S (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14903__A1 (.I(_06859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14906__A1 (.I(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14908__I (.I(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14909__I1 (.I(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14915__I (.I(_06786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14916__A1 (.I(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14921__B2 (.I(_06859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14923__A1 (.I(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14924__A2 (.I(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14928__A1 (.I(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14931__A1 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14939__A1 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14939__B (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14942__A1 (.I(\filters.band[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14942__A2 (.I(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14947__A1 (.I(_06747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14948__A1 (.I(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14949__A1 (.I(\filters.band[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14949__B (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14951__A1 (.I(_06745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14952__A1 (.I(_06745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14954__I1 (.I(\filters.band[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14955__A1 (.I(_06793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14956__A1 (.I(\filters.band[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14956__B (.I(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14958__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14958__A2 (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14961__I (.I(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14962__I (.I(\filters.low[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14965__A2 (.I(_06936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14965__B (.I(_06937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14967__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14967__A2 (.I(_06939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14968__I (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14969__A2 (.I(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14969__C (.I(_06941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14974__A3 (.I(\channels.sample1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14974__A4 (.I(\channels.sample2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14975__A2 (.I(\channels.sample1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14975__B1 (.I(\channels.sample2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14977__A2 (.I(\channels.sample3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14978__A1 (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14980__A2 (.I(_06936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14981__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14981__A2 (.I(_06939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14982__A1 (.I(_06945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14983__B (.I(_06945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14984__A1 (.I(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14985__A1 (.I(\filters.high[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14985__A2 (.I(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14986__A1 (.I(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14990__A1 (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14990__A2 (.I(\channels.sample3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14991__A1 (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14993__A3 (.I(\channels.sample1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14993__A4 (.I(\channels.sample2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14994__A2 (.I(\channels.sample1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14994__B1 (.I(\channels.sample2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14996__A2 (.I(\channels.sample3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15002__A2 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15003__A2 (.I(_06973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15004__A1 (.I(_06959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15004__A2 (.I(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15006__A1 (.I(_06959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15006__A2 (.I(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15006__B (.I(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15007__A1 (.I(\filters.high[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15007__A2 (.I(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15008__A1 (.I(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15009__I (.I(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15010__A1 (.I(\filters.high[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15010__A2 (.I(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15011__A2 (.I(_06973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15012__A1 (.I(_06959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15012__A2 (.I(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15016__A1 (.I(\filters.filt_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15016__A2 (.I(\filters.filt_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15016__A3 (.I(\channels.sample1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15016__A4 (.I(\channels.sample2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15017__A1 (.I(\filters.filt_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15017__A2 (.I(\channels.sample1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15017__B1 (.I(\channels.sample2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15017__B2 (.I(\filters.filt_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15019__A1 (.I(\filters.filt_3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15019__A2 (.I(\channels.sample3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15024__A2 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15026__A2 (.I(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15027__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15030__B (.I(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15032__B (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15033__A2 (.I(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15034__A1 (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15034__A2 (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15036__I (.I(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15040__A1 (.I(\filters.filt_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15040__A2 (.I(\filters.filt_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15040__A3 (.I(\channels.sample1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15040__A4 (.I(\channels.sample2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15041__A2 (.I(\channels.sample1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15041__B1 (.I(\channels.sample2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15043__A2 (.I(\channels.sample3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15050__A1 (.I(\filters.low[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15052__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15058__A1 (.I(_07005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15059__B (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15062__A1 (.I(_05994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15063__A1 (.I(_05994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15072__A2 (.I(\channels.sample3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15073__A2 (.I(\channels.sample2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15074__A2 (.I(\channels.sample1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15079__A1 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15085__B (.I(_07052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15088__A1 (.I(\filters.high[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15088__A2 (.I(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15088__B (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15089__A1 (.I(_07054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15091__I (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15101__A2 (.I(\channels.sample2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15102__A2 (.I(\channels.sample1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15109__A3 (.I(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15112__A1 (.I(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15113__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15118__I (.I(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15119__I (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15120__A1 (.I(\filters.high[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15120__A2 (.I(_07085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15120__B (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15121__A1 (.I(_07058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15121__A2 (.I(_07084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15122__I (.I(_06937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15123__A1 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15123__A2 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15128__A2 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15131__A2 (.I(\channels.sample3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15132__A2 (.I(\channels.sample2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15133__A2 (.I(\channels.sample1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15136__A2 (.I(_07101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15138__A1 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15145__B (.I(_07110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15147__A2 (.I(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15147__C (.I(_06773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15165__A2 (.I(\channels.sample2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15166__A2 (.I(\channels.sample1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15173__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15173__A2 (.I(_07101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15178__A1 (.I(_06937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15178__A2 (.I(_07142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15179__A2 (.I(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15179__C (.I(_06773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15180__A1 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15180__A2 (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15185__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15188__A2 (.I(\channels.sample3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15189__A2 (.I(\channels.sample2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15190__A2 (.I(\channels.sample1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15196__A1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15201__B (.I(_07110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15203__A1 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15203__A2 (.I(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15203__C (.I(_06773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15218__A2 (.I(\channels.sample2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15219__A2 (.I(\channels.sample1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15223__A2 (.I(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15223__A3 (.I(_07185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15227__A1 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15229__A2 (.I(_07191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15230__A1 (.I(_07169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15230__A2 (.I(_07172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15231__A2 (.I(_07169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15231__A3 (.I(_07172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15232__A1 (.I(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15233__A1 (.I(\filters.high[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15233__A2 (.I(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15234__A1 (.I(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15235__A1 (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15235__A2 (.I(_07185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15236__A1 (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15236__A2 (.I(_07185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15241__A2 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15244__A2 (.I(\channels.sample3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15245__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15245__A2 (.I(\channels.sample2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15246__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15246__A2 (.I(\channels.sample1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15249__A2 (.I(_07210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15250__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15250__A2 (.I(_07210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15254__A2 (.I(_07191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15255__B (.I(_07110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15257__I (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15258__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15258__A2 (.I(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15258__C (.I(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15260__A1 (.I(_07169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15260__A2 (.I(_07172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15261__A2 (.I(_07191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15274__A2 (.I(\channels.sample3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15275__A2 (.I(\channels.sample2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15276__A2 (.I(\channels.sample1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15280__A2 (.I(_07240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15281__A2 (.I(_07240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15286__A1 (.I(\filters.high[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15286__A2 (.I(_07085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15286__B (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15287__A1 (.I(_07058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15287__A2 (.I(_07246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15289__A2 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15294__A1 (.I(_07250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15294__A2 (.I(_07253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15297__A1 (.I(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15297__A2 (.I(_05878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15303__B (.I(_07052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15305__A2 (.I(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15305__B (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15307__A1 (.I(_07250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15307__A2 (.I(_07253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15309__A1 (.I(_05993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15312__A1 (.I(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15320__B (.I(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15322__A1 (.I(\filters.high[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15322__A2 (.I(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15323__A1 (.I(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15324__A2 (.I(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15325__A1 (.I(_05993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15326__A1 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15331__B (.I(_07110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15333__A2 (.I(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15333__C (.I(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15342__A2 (.I(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15343__A1 (.I(\filters.low[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15344__A1 (.I(_07299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15345__A1 (.I(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15346__A2 (.I(_07085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15346__B (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15347__A1 (.I(_07058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15348__A1 (.I(\filters.low[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15349__A1 (.I(\filters.low[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15350__A1 (.I(_07299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15351__A1 (.I(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15353__A1 (.I(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15355__A2 (.I(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15355__B (.I(_07310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15357__A2 (.I(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15358__A1 (.I(\filters.low[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15359__A2 (.I(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15362__I (.I(\filters.low[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15363__A1 (.I(_07317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15367__A1 (.I(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15369__A1 (.I(_07005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15370__B (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15371__A2 (.I(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15374__A1 (.I(_07317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15375__A1 (.I(_07317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15378__I (.I(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15379__B (.I(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15380__A1 (.I(_07058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15381__I (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15382__A2 (.I(_06522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15383__A2 (.I(_06625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15390__B2 (.I(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15392__I (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15399__A2 (.I(_06625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15404__A2 (.I(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15406__A1 (.I(\filters.low[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15409__A2 (.I(_06860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15416__A1 (.I(_07085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15417__I (.I(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15418__B (.I(_07368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15421__A1 (.I(\filters.low[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15421__A2 (.I(_06860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15437__A2 (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15439__I (.I(\filters.high[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15441__B (.I(_07380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15448__A1 (.I(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15451__A1 (.I(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15452__A2 (.I(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15452__C (.I(_06941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15456__A2 (.I(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15457__I0 (.I(_07401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15460__A1 (.I(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15464__A1 (.I(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15465__A2 (.I(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15469__A1 (.I(_07401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15469__A2 (.I(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15470__I0 (.I(_07413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15471__A1 (.I(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15473__B (.I(_07052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15475__A2 (.I(_07005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15475__B (.I(_07310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15479__A1 (.I(_07401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15480__A1 (.I(_07413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15481__B2 (.I(_07380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15482__A1 (.I(_07413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15483__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15487__I (.I(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15488__A2 (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15488__B (.I(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15489__A1 (.I(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15489__A2 (.I(_07431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15492__A1 (.I(_07435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15492__A2 (.I(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15496__B (.I(_07052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15498__A2 (.I(_07005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15498__B (.I(_07310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15500__A2 (.I(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15502__A1 (.I(_07435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15506__A1 (.I(_07435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15507__A1 (.I(_07435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15509__B (.I(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15511__B (.I(_07368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15518__B (.I(_06937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15519__A2 (.I(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15519__C (.I(_06941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15520__I (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15521__A1 (.I(\filters.mode_vol[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15521__A2 (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15521__C (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15522__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15522__B1 (.I(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15522__B2 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15523__C (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15524__I (.I(_07464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15526__A1 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15526__A2 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15526__B (.I(_07464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15529__A1 (.I(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15529__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15529__A3 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15531__A1 (.I(\channels.sample3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15532__A1 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15533__A1 (.I(\channels.sample2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15534__A1 (.I(\channels.sample1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15536__A2 (.I(_07476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15537__A2 (.I(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15539__I (.I(_07464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15540__A2 (.I(_07476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15542__A1 (.I(\channels.sample3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15544__A1 (.I(\channels.sample2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15545__A1 (.I(\channels.sample1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15547__A2 (.I(_07486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15551__A2 (.I(_07486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15553__A1 (.I(\channels.sample3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15555__A1 (.I(\channels.sample2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15555__A2 (.I(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15556__A1 (.I(\channels.sample1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15558__A2 (.I(_07496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15564__I (.I(_07464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15565__A1 (.I(\filters.sample_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15567__A2 (.I(_07496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15569__A1 (.I(\channels.sample3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15570__C (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15571__A1 (.I(\channels.sample2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15572__A1 (.I(\channels.sample1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15574__A1 (.I(\filters.sample_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15574__A2 (.I(_07511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15578__B (.I(_07368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15580__A1 (.I(\filters.sample_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15580__A2 (.I(_07511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15581__A1 (.I(\channels.sample3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15583__A1 (.I(\channels.sample2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15583__A2 (.I(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15584__A1 (.I(\channels.sample1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15586__A2 (.I(_07522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15592__A1 (.I(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15594__A2 (.I(_07522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15596__A1 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15597__C (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15598__A1 (.I(\channels.sample2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15598__A2 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15599__A1 (.I(\channels.sample1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15601__A2 (.I(_07536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15605__B (.I(_07368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15607__A2 (.I(_07536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15608__A1 (.I(\channels.sample3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15609__C (.I(_06202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15610__A1 (.I(\channels.sample2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15610__A2 (.I(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15611__A1 (.I(\channels.sample1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15613__A2 (.I(_07547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15619__A1 (.I(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15621__A2 (.I(_07547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15623__A1 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15624__C (.I(_06733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15625__A1 (.I(\channels.sample2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15626__A1 (.I(\channels.sample1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15628__A2 (.I(_07561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15632__I (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15633__I (.I(_07566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15635__A2 (.I(_07561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15637__A1 (.I(\channels.sample3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15639__A1 (.I(\channels.sample2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15640__A1 (.I(\channels.sample1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15642__A2 (.I(_07574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15648__A1 (.I(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15649__A2 (.I(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15650__A2 (.I(_07574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15652__A1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15654__A1 (.I(\channels.sample2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15655__A1 (.I(\channels.sample1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15657__A2 (.I(_07588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15662__A2 (.I(_07588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15663__A1 (.I(\channels.sample3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15665__A1 (.I(\channels.sample2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15666__A1 (.I(\channels.sample1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15668__A2 (.I(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15674__A1 (.I(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15675__A1 (.I(\filters.sample_buff[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15675__A2 (.I(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15676__A2 (.I(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15677__A1 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15679__A1 (.I(\channels.sample2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15680__A1 (.I(\channels.sample1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15682__A1 (.I(\filters.sample_buff[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15682__A2 (.I(_07611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15687__I (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15689__A1 (.I(\filters.sample_buff[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15689__A2 (.I(_07611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15691__A1 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15693__A1 (.I(\filters.sample_buff[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15694__B (.I(\filters.sample_buff[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15697__A1 (.I(\filters.sample_buff[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15698__A1 (.I(_07617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15699__A1 (.I(\filters.sample_buff[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15699__A2 (.I(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15702__A1 (.I(\filters.sample_buff[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15707__I (.I(\filters.sample_buff[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15708__A1 (.I(\filters.sample_buff[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15715__C (.I(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15726__A2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15729__I (.I(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15731__I (.I(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15732__A1 (.I(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15732__B (.I(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15733__A2 (.I(_07651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15734__A2 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15734__A3 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15735__I (.I(_07654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15736__I (.I(_07655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15739__I (.I(_07658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15740__A1 (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15740__A2 (.I(_07659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15740__B (.I(_07310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15743__I (.I(_07658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15744__I (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15745__I (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15746__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15747__A1 (.I(_07661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15749__A1 (.I(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15751__A1 (.I(_05994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15751__B (.I(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15752__A2 (.I(_07651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15754__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15755__A1 (.I(_07669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15756__I (.I(_07655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15758__A1 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15759__A1 (.I(_07672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15761__I (.I(_07658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15762__I (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15763__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15766__A1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15769__A1 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15771__I (.I(_07654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15772__I (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15774__A1 (.I(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15776__A1 (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15776__B (.I(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15777__A2 (.I(_07651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15778__I (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15779__I (.I(_07687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15780__B (.I(_07688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15781__A2 (.I(_07651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15783__I (.I(_07658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15784__I (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15788__A1 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15793__I (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15794__A2 (.I(_07698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15795__A1 (.I(\filters.low[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15797__A1 (.I(_07317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15797__B (.I(_07688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15798__A2 (.I(_07659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15799__A2 (.I(_07698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15800__I (.I(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15801__I (.I(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15804__A2 (.I(_07698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15807__A2 (.I(_07698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15810__I (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15815__I (.I(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15816__I (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15817__I (.I(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15818__A1 (.I(\filters.low[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15820__I (.I(_07655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15821__I (.I(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15823__A2 (.I(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15823__C (.I(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15824__B (.I(_07688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15825__A2 (.I(_07659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15827__A1 (.I(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15830__A1 (.I(_07401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15833__A1 (.I(_07413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15836__I (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15837__A2 (.I(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15837__C (.I(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15839__A2 (.I(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15839__C (.I(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15840__A2 (.I(_07655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15841__A2 (.I(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15841__C (.I(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15842__B (.I(_07688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15843__A2 (.I(_07659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15844__I (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15845__A1 (.I(_07733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15846__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15846__A2 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15847__A3 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15848__A1 (.I(_07733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15849__A1 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15851__A1 (.I(_07617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15857__I (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15858__A2 (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15858__A3 (.I(_07743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15859__I (.I(_07566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15864__A2 (.I(_07748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15867__A1 (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15867__A2 (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15870__A1 (.I(_07617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15874__A1 (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15875__A1 (.I(_07733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15881__I (.I(_07762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15884__A1 (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15884__A2 (.I(_07764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15884__C (.I(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15905__I (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15915__A2 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15959__A2 (.I(_07839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15962__A2 (.I(_07839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15974__I (.I(_07748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15978__A1 (.I(_07617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15979__I (.I(_07743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16012__I (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16013__B1 (.I(_07891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16014__A1 (.I(_07859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16052__A2 (.I(_07839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16057__A2 (.I(_07924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16065__A1 (.I(_07859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16086__A1 (.I(_07950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16086__A2 (.I(_07959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16087__A1 (.I(_07924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16088__A1 (.I(_07924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16092__B (.I(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16093__A2 (.I(_07748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16095__A2 (.I(_07945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16096__A1 (.I(_07944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16113__A1 (.I(_07977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16113__A3 (.I(_07989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16114__A1 (.I(_07959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16115__A1 (.I(_07959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16116__A1 (.I(_07950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16119__A1 (.I(_07859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16123__I (.I(_07977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16124__A2 (.I(_07989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16125__A2 (.I(_07989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16150__A1 (.I(_07764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16176__C (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16177__A1 (.I(_07764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16201__C (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16202__A1 (.I(_07764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16223__B1 (.I(_07891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16223__C (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16244__A1 (.I(_07748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16247__I (.I(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16248__A2 (.I(_07945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16248__B (.I(_08119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16257__B (.I(_07762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16260__A2 (.I(_07891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16260__B (.I(_08119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16263__A2 (.I(_07743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16264__I (.I(_07687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16265__A2 (.I(_07891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16265__B (.I(_08134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16266__A1 (.I(_07945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16267__A1 (.I(\filters.sample_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16267__A2 (.I(_07743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16268__A1 (.I(_07944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16269__I (.I(_07762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16273__A1 (.I(_07944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16276__A1 (.I(_07944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16283__I (.I(_07762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16293__A1 (.I(\filters.sample_buff[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16295__A1 (.I(\filters.sample_buff[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16297__A1 (.I(\filters.sample_buff[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16299__I (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16300__I (.I(_08157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16301__A1 (.I(\filters.sample_buff[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16303__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16306__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16309__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16309__A2 (.I(_07859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16311__A1 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16342__A1 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16344__A1 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16344__A2 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16344__B (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16357__A1 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16361__A1 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16364__B1 (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16366__B1 (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16368__A2 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16368__B1 (.I(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16370__A2 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16370__B1 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16372__A2 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16372__B1 (.I(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16374__A1 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16376__A1 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16376__A2 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16376__B (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16378__A1 (.I(\channels.ch3_env[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16380__A1 (.I(\channels.ch3_env[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16382__A1 (.I(\channels.ch3_env[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16384__A1 (.I(\channels.ch3_env[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16388__A1 (.I(\channels.ch3_env[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16389__A1 (.I(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16390__A1 (.I(\channels.ch3_env[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16392__A1 (.I(\channels.ch3_env[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16393__A1 (.I(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16394__A1 (.I(\channels.ch3_env[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16398__I (.I(_08213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16399__A2 (.I(_08213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16400__A2 (.I(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16401__I (.I(_08216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16405__I (.I(_08219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16409__I (.I(_08213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16420__I (.I(_08219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16422__I (.I(_08216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16424__I (.I(_08213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16435__I (.I(_08219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16437__I (.I(_08216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16450__A2 (.I(_08219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16452__A1 (.I(\tt_um_rejunity_sn76489.control_noise[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16453__A1 (.I(_07839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16459__I (.I(_08259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16460__A2 (.I(_08260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16464__I (.I(_08263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16467__A2 (.I(_08266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16469__A1 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16471__B (.I(_08119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16474__B (.I(_08119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16477__I (.I(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16478__B (.I(_08274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16480__B (.I(_08134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16485__A2 (.I(_07945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16486__I (.I(_08263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16490__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16492__I (.I(_08259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16493__A2 (.I(_08285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16494__I (.I(_07566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16495__B (.I(_08287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16496__I (.I(_08157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16498__I (.I(_08263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16502__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16502__A2 (.I(_08290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16506__I (.I(_08259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16507__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16508__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16511__A1 (.I(_08297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16512__I (.I(_08263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16515__A2 (.I(_08305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16515__B (.I(_08274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16517__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16519__B (.I(_08266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16521__A2 (.I(_08305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16521__B (.I(_08274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16527__B (.I(_08315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16528__A2 (.I(_08312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16532__B (.I(_08315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16533__A2 (.I(_08312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16539__A2 (.I(_08312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16544__A1 (.I(_08297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16545__A2 (.I(_08305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16545__B (.I(_08274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16549__A1 (.I(_08260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16550__A2 (.I(_08285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16551__B (.I(_08287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16552__I (.I(_08157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16554__A2 (.I(_08337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16556__A1 (.I(_08336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16557__A2 (.I(_08337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16557__B (.I(_08134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16558__A2 (.I(_08337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16562__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16564__A2 (.I(_08285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16565__B (.I(_08287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16570__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16570__A2 (.I(_08290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16573__A1 (.I(_08336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16574__I (.I(_08259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16575__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16576__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16579__A1 (.I(_08354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16580__I (.I(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16581__A2 (.I(_08305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16581__B (.I(_08360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16583__A1 (.I(\tt_um_rejunity_sn76489.control_tone_freq[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16585__B (.I(_08315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16588__B (.I(_08360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16594__A2 (.I(_08368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16595__A1 (.I(_08336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16599__A2 (.I(_08368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16600__A1 (.I(_08336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16601__I (.I(_08157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16605__A2 (.I(_08368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16606__A1 (.I(_08377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16610__A1 (.I(_08354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16611__B (.I(_08360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16615__A1 (.I(_08260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16616__A2 (.I(_08297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16617__B (.I(_08287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16619__A2 (.I(_08391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16621__A1 (.I(_08377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16622__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16622__A2 (.I(_08391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16622__B (.I(_08134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16623__A1 (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16623__A2 (.I(_08391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16624__A1 (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16625__I (.I(_08395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16627__A1 (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16627__A2 (.I(_08395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16630__B1 (.I(_08400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16631__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16631__B1 (.I(_08400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16632__B1 (.I(_08400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16633__A1 (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16633__B1 (.I(_08400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16634__I (.I(_08395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16635__I (.I(_08401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16637__I (.I(_08403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16640__A1 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16642__I (.I(_08401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16643__I (.I(_08403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16646__A1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16648__I (.I(_08401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16649__I (.I(_08403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16650__A1 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16653__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16654__I (.I(_08401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16655__I (.I(_08403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16658__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16659__A1 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16660__A1 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16661__A1 (.I(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16668__A1 (.I(_08290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16669__A2 (.I(_08285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16670__I (.I(_07566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16671__B (.I(_08418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16676__A2 (.I(_08290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16679__A1 (.I(_08377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16684__A1 (.I(_08354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16685__B (.I(_08360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16689__B (.I(_08315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16691__B (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16696__A2 (.I(_08368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16697__A1 (.I(_08377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16698__I (.I(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16702__A2 (.I(_08266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16703__A1 (.I(_08441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16707__A2 (.I(_08266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16708__A1 (.I(_08441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16712__A1 (.I(_08354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16713__A2 (.I(_08312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16713__B (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16717__A1 (.I(_08260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16718__A2 (.I(_08297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16719__B (.I(_08418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16721__A2 (.I(_08459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16723__A1 (.I(_08441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16724__I (.I(_07687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16725__A2 (.I(_08459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16726__A2 (.I(_08459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16728__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16728__A3 (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16729__A2 (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16735__A1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16736__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16738__A1 (.I(_08472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16739__I (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16741__A1 (.I(_08474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16742__I (.I(_07687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16744__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16747__A1 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16748__B (.I(_08418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16750__A1 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16752__A2 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16753__A3 (.I(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16759__A1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16761__A1 (.I(_08472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16763__B (.I(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16764__A1 (.I(_08474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16766__B (.I(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16767__A1 (.I(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16770__A1 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16771__B (.I(_08418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16772__B (.I(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16773__A1 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16778__B (.I(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16779__A1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16782__A1 (.I(_08472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16784__A1 (.I(_08474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16786__A1 (.I(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16789__A1 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16790__B (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16792__A1 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16801__I (.I(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16802__I (.I(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16803__A1 (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16804__I (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16806__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16808__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16810__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16813__A1 (.I(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16816__I (.I(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16817__I (.I(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16818__A1 (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16819__I (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16822__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16824__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16826__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16828__A2 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16830__I (.I(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16831__I (.I(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16833__I (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16834__A1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16836__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16838__A1 (.I(_08474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16840__A1 (.I(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16841__B2 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16843__I (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16844__I (.I(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16846__I (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16847__A1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16849__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16851__A1 (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16853__A1 (.I(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16855__A2 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16856__A1 (.I(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16856__B (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16860__A1 (.I(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16860__B (.I(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16863__C (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16864__C (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16866__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16866__B (.I(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16867__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16868__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16869__A3 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16870__A1 (.I(_06941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16872__B (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16874__B (.I(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16878__A1 (.I(_08441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16879__A1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16879__A2 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16879__B (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16880__I (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16881__I (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16882__A2 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16882__C (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16883__A1 (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16884__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16884__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16885__A2 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16885__A3 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16887__A1 (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16887__A3 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16887__A4 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16895__A2 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16895__B (.I(\channels.clk_div[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16896__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16896__A2 (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16896__A3 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16896__A4 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16899__A1 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16899__A2 (.I(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16904__B (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16908__A1 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16909__A1 (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16911__I0 (.I(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16911__S (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16921__A1 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16921__A2 (.I(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16922__I (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16923__S (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16925__S (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16927__I0 (.I(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16927__S (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16929__S (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16931__S (.I(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16943__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16943__A2 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16943__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16944__I (.I(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16945__S (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16947__S (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16949__I0 (.I(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16949__S (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16951__S (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16953__S (.I(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16955__A1 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16956__A2 (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16956__B (.I(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16957__A1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16957__A2 (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16958__A2 (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16958__B (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16959__A1 (.I(_08472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16959__A2 (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16960__A1 (.I(\tt_um_rejunity_sn76489.control_noise[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16960__A2 (.I(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16961__A1 (.I(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16961__A2 (.I(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16961__C (.I(_07733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17002__CLK (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17009__CLK (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17058__D (.I(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17085__D (.I(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17086__D (.I(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17087__D (.I(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17094__CLK (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17108__CLK (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17238__CLK (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17274__CLK (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17279__CLK (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17326__CLK (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17378__CLK (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17447__CLK (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17512__D (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17513__D (.I(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17514__D (.I(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17515__D (.I(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17531__CLK (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17535__CLK (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17576__D (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17577__D (.I(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17578__D (.I(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17579__D (.I(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17593__CLK (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17598__CLK (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17602__CLK (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17602__D (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17603__D (.I(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17604__D (.I(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17637__D (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17673__CLK (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17697__D (.I(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17767__CLK (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17775__CLK (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_0__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_10__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_11__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_12__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_13__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_14__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_15__f_clk_I (.I(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_16__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_17__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_18__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_19__f_clk_I (.I(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_1__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_20__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_21__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_22__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_23__f_clk_I (.I(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_24__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_25__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_26__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_27__f_clk_I (.I(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_28__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_29__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_2__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_30__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_31__f_clk_I (.I(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_3__f_clk_I (.I(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_4__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_5__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_6__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_7__f_clk_I (.I(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_8__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_5_9__f_clk_I (.I(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_clk_I (.I(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_126_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_128_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_129_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_130_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_131_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_132_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_133_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_134_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_135_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_136_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_138_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_139_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_140_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_141_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_142_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_143_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_144_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_145_clk_I (.I(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_146_clk_I (.I(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_147_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_148_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_149_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_150_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_151_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_152_clk_I (.I(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_153_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_154_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_155_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_156_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_157_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_158_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_159_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_160_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_161_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_162_clk_I (.I(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_163_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_164_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_165_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_166_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_167_clk_I (.I(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_168_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_169_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_170_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_171_clk_I (.I(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_172_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_173_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_174_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_175_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_176_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_177_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_178_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_179_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_180_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_181_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_183_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_184_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_185_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_186_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_187_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_188_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_190_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_191_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_192_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_193_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_194_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_195_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_196_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_197_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_199_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clk_I (.I(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_200_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_201_clk_I (.I(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_202_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_203_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_204_clk_I (.I(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_205_clk_I (.I(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_207_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_208_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_209_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_210_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_211_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_212_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_213_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_214_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_215_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_216_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_217_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_218_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_219_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_220_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_221_clk_I (.I(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_222_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_223_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_224_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_225_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_226_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_227_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_228_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_229_clk_I (.I(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_230_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_231_clk_I (.I(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_232_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_233_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_234_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_235_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_236_clk_I (.I(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_237_clk_I (.I(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_238_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_239_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_240_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_241_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_242_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_243_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_244_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_245_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_246_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clk_I (.I(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clk_I (.I(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clk_I (.I(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clk_I (.I(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_clk_I (.I(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clk_I (.I(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_clk_I (.I(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clk_I (.I(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_clk_I (.I(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_clk_I (.I(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_clk_I (.I(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_clk_I (.I(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_clk_I (.I(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_clk_I (.I(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_clk_I (.I(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clk_I (.I(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(bus_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(bus_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(bus_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(bus_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(bus_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(bus_we));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(bus_cyc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(bus_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(bus_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(bus_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer13_I (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer14_I (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer1_I (.I(_07380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer20_I (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer25_I (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer31_I (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer35_I (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer3_I (.I(_06859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer42_I (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer43_I (.I(_07380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer5_I (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer6_I (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer8_I (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_179_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Left_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Left_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Left_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Left_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Left_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Left_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Left_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Left_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Left_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Left_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Left_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Left_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Left_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Left_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Left_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Left_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Left_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Left_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Left_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Left_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Left_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Left_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Left_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Left_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Left_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Left_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Left_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Left_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Left_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Left_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Left_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Left_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Left_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Left_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Left_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Left_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Left_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Left_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_569 ();
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08482_ (.I(net5),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08483_ (.I(net4),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08484_ (.A1(_01012_),
    .A2(net3),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08485_ (.A1(net2),
    .A2(net1),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08486_ (.A1(_01011_),
    .A2(_01013_),
    .A3(_01014_),
    .ZN(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _08487_ (.A1(net6),
    .A2(net15),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08488_ (.A1(_01015_),
    .A2(_01016_),
    .ZN(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08489_ (.A1(\filters.res_filt[5] ),
    .A2(_01017_),
    .ZN(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08490_ (.A1(_01015_),
    .A2(_01016_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08491_ (.I(_01019_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08492_ (.A1(net12),
    .A2(_01020_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08493_ (.A1(_01018_),
    .A2(_01021_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08494_ (.I(net16),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08495_ (.A1(net13),
    .A2(_01017_),
    .ZN(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08496_ (.A1(\filters.res_filt[6] ),
    .A2(_01019_),
    .ZN(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08497_ (.A1(_01023_),
    .A2(_01024_),
    .A3(_01025_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08498_ (.I(_01026_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08499_ (.I(_01023_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08500_ (.I(net11),
    .ZN(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08501_ (.A1(_01029_),
    .A2(_01019_),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08502_ (.A1(\filters.res_filt[4] ),
    .A2(_01020_),
    .B(_01030_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08503_ (.A1(_01028_),
    .A2(_01031_),
    .ZN(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08504_ (.I(_01032_),
    .Z(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08505_ (.A1(_01022_),
    .A2(_01027_),
    .A3(_00129_),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08506_ (.I(_01026_),
    .ZN(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08507_ (.A1(net14),
    .A2(_01017_),
    .ZN(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08508_ (.A1(\filters.res_filt[7] ),
    .A2(_01019_),
    .ZN(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _08509_ (.A1(_01028_),
    .A2(_01035_),
    .A3(_01036_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08510_ (.I(_01037_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08511_ (.A1(_01034_),
    .A2(_01031_),
    .B(_01038_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08512_ (.I(_01034_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08513_ (.I(_01023_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08514_ (.A1(_01040_),
    .A2(_01022_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08515_ (.I(net12),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08516_ (.A1(_01042_),
    .A2(_01017_),
    .B(_01018_),
    .ZN(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08517_ (.A1(_01043_),
    .A2(_01032_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08518_ (.A1(_01032_),
    .A2(_01041_),
    .B(_01044_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08519_ (.A1(_00131_),
    .A2(_01045_),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08520_ (.I(_01044_),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08521_ (.I(_01037_),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08522_ (.A1(_01027_),
    .A2(_01047_),
    .B(_01048_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08523_ (.A1(_01033_),
    .A2(_01039_),
    .B1(_01046_),
    .B2(_01049_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08524_ (.A1(_01043_),
    .A2(_01026_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08525_ (.A1(_00129_),
    .A2(_01050_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08526_ (.I(_01040_),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08527_ (.A1(_01052_),
    .A2(_01022_),
    .B(_01026_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08528_ (.A1(_01039_),
    .A2(_01053_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08529_ (.A1(_01051_),
    .A2(_01054_),
    .Z(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08530_ (.I(_01055_),
    .Z(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08531_ (.A1(_01027_),
    .A2(_00129_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08532_ (.A1(_01056_),
    .A2(_01046_),
    .B(_01038_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08533_ (.A1(_01056_),
    .A2(_01046_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08534_ (.A1(_00131_),
    .A2(_01031_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08535_ (.A1(_01059_),
    .A2(_01047_),
    .B(_01038_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08536_ (.A1(_01058_),
    .A2(_01060_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08537_ (.A1(_01057_),
    .A2(_01061_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08538_ (.I(_01041_),
    .Z(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08539_ (.A1(_01059_),
    .A2(_01044_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08540_ (.A1(_01048_),
    .A2(_00130_),
    .B(_01062_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08541_ (.A1(_01060_),
    .A2(_01063_),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08542_ (.I(_01064_),
    .Z(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08543_ (.I(_01038_),
    .Z(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08544_ (.A1(_01027_),
    .A2(_00130_),
    .B(_01050_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08545_ (.A1(_01056_),
    .A2(_00132_),
    .A3(_01065_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08546_ (.A1(_00131_),
    .A2(_01048_),
    .A3(_01047_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08547_ (.A1(_01066_),
    .A2(_01067_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08548_ (.A1(_01047_),
    .A2(_01053_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08549_ (.I0(_01031_),
    .I1(_01068_),
    .S(_01037_),
    .Z(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08550_ (.I(_01069_),
    .Z(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08551_ (.A1(_01022_),
    .A2(_01048_),
    .B(_01054_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08552_ (.A1(_00132_),
    .A2(_01065_),
    .B(_01057_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08553_ (.A1(_01032_),
    .A2(_00130_),
    .B(_01034_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08554_ (.A1(_00132_),
    .A2(_01070_),
    .B(_01053_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08555_ (.I(_01023_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08556_ (.I(\clk_ctr[0] ),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08557_ (.A1(\clk_trg[0] ),
    .A2(_01072_),
    .B(\clk_ctr[1] ),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08558_ (.A1(\clk_trg[1] ),
    .A2(_01073_),
    .ZN(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08559_ (.I(\clk_trg[0] ),
    .ZN(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08560_ (.I(\clk_trg[1] ),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08561_ (.A1(_01076_),
    .A2(\clk_ctr[1] ),
    .B(_01072_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08562_ (.A1(_01075_),
    .A2(_01077_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08563_ (.A1(_01074_),
    .A2(_01078_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08564_ (.A1(_01071_),
    .A2(_01079_),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08565_ (.A1(\channels.clk_div[0] ),
    .A2(_01080_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08566_ (.I(\channels.clk_div[2] ),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08567_ (.I(\channels.clk_div[1] ),
    .Z(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08568_ (.A1(_01082_),
    .A2(_01083_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08569_ (.I(_01084_),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08570_ (.I(_01085_),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08571_ (.I(_01086_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08572_ (.I(_01087_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08573_ (.I(_01088_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08574_ (.I(_01089_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08575_ (.I(_01090_),
    .Z(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08576_ (.I(_01091_),
    .Z(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08577_ (.I(_01092_),
    .Z(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08578_ (.A1(_01081_),
    .A2(_01093_),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08579_ (.I(_01094_),
    .Z(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08580_ (.I0(\channels.accum[0][23] ),
    .I1(\channels.accum[1][23] ),
    .I2(\channels.accum[2][23] ),
    .I3(\channels.accum[3][23] ),
    .S0(_00009_),
    .S1(_00010_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08581_ (.I(_01096_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08582_ (.I(_01028_),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08583_ (.A1(_01098_),
    .A2(_01094_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08584_ (.I(_01099_),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08585_ (.I(_01100_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08586_ (.A1(_01095_),
    .A2(_01097_),
    .B1(_01101_),
    .B2(\channels.ring_outs[2] ),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08587_ (.I(_01102_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08588_ (.I(\channels.clk_div[0] ),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08589_ (.A1(_01074_),
    .A2(_01078_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08590_ (.A1(net16),
    .A2(_01104_),
    .ZN(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08591_ (.A1(_01103_),
    .A2(_01105_),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08592_ (.I(_01082_),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08593_ (.I(_01107_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08594_ (.I(_01083_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08595_ (.A1(_01108_),
    .A2(_01109_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08596_ (.A1(_01106_),
    .A2(_01110_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08597_ (.I(_01111_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08598_ (.A1(_01098_),
    .A2(_01111_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08599_ (.I(_01113_),
    .Z(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08600_ (.I(_01114_),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08601_ (.A1(_01097_),
    .A2(_01112_),
    .B1(_01115_),
    .B2(\channels.ring_outs[1] ),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08602_ (.I(_01116_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08603_ (.I(\channels.lfsr[3][0] ),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08604_ (.I(_01117_),
    .Z(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08605_ (.I(\channels.lfsr[3][1] ),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08606_ (.I(_01118_),
    .Z(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08607_ (.I(\channels.lfsr[3][2] ),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08608_ (.I(_01119_),
    .Z(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08609_ (.I(\channels.lfsr[3][3] ),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08610_ (.I(_01120_),
    .Z(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08611_ (.I(\channels.lfsr[3][4] ),
    .Z(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08612_ (.I(_01121_),
    .Z(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08613_ (.I(\channels.lfsr[3][5] ),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08614_ (.I(_01122_),
    .Z(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08615_ (.I(\channels.lfsr[3][6] ),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08616_ (.I(_01123_),
    .Z(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08617_ (.I(\channels.lfsr[3][7] ),
    .Z(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08618_ (.I(_01124_),
    .Z(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08619_ (.I(\channels.lfsr[3][8] ),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08620_ (.I(_01125_),
    .Z(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08621_ (.I(\channels.lfsr[3][9] ),
    .Z(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08622_ (.I(_01126_),
    .Z(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08623_ (.I(\channels.lfsr[3][10] ),
    .Z(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08624_ (.I(_01127_),
    .Z(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08625_ (.I(\channels.lfsr[3][11] ),
    .Z(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08626_ (.I(_01128_),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08627_ (.I(\channels.lfsr[3][12] ),
    .Z(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08628_ (.I(_01129_),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08629_ (.I(\channels.lfsr[3][13] ),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08630_ (.I(_01130_),
    .Z(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08631_ (.I(\channels.lfsr[3][14] ),
    .Z(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08632_ (.I(_01131_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08633_ (.I(\channels.lfsr[3][15] ),
    .Z(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08634_ (.I(_01132_),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08635_ (.I(\channels.lfsr[3][16] ),
    .Z(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08636_ (.I(_01133_),
    .Z(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08637_ (.I(\channels.lfsr[3][17] ),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08638_ (.I(_01134_),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08639_ (.I(\channels.lfsr[3][18] ),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08640_ (.I(_01135_),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08641_ (.I(\channels.lfsr[3][19] ),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08642_ (.I(_01136_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08643_ (.I(\channels.lfsr[3][20] ),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08644_ (.I(_01137_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08645_ (.I(\channels.lfsr[3][21] ),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08646_ (.I(_01138_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08647_ (.I(\channels.lfsr[3][22] ),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08648_ (.I(_01139_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08649_ (.I(\channels.env_vol[3][0] ),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08650_ (.I(_01140_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08651_ (.I(\channels.env_vol[3][1] ),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08652_ (.I(_01141_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08653_ (.I(\channels.env_vol[3][2] ),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08654_ (.I(_01142_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08655_ (.I(\channels.env_vol[3][3] ),
    .Z(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08656_ (.I(_01143_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08657_ (.I(\channels.env_vol[3][4] ),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08658_ (.I(_01144_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08659_ (.I(\channels.env_vol[3][5] ),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08660_ (.I(_01145_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08661_ (.I(\channels.env_vol[3][6] ),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08662_ (.I(_01146_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08663_ (.I(\channels.env_vol[3][7] ),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08664_ (.I(_01147_),
    .Z(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08665_ (.I(_00009_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08666_ (.I(_01148_),
    .Z(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08667_ (.I(_01149_),
    .Z(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08668_ (.I(_01150_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08669_ (.I(_01151_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08670_ (.I(_01152_),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08671_ (.I(_01153_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08672_ (.I(_01154_),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08673_ (.I(_01155_),
    .Z(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08674_ (.I(_01156_),
    .Z(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08675_ (.I(_01157_),
    .Z(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08676_ (.I(_01158_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08677_ (.I(_01159_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08678_ (.I(_01160_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08679_ (.I(_01161_),
    .Z(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08680_ (.I(_00010_),
    .Z(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08681_ (.I(_01163_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08682_ (.I(_01164_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08683_ (.I(_01165_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08684_ (.I(_01166_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08685_ (.I(_01167_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08686_ (.I(_01168_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08687_ (.I(_01169_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08688_ (.I(_01170_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08689_ (.I(_01171_),
    .Z(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08690_ (.I(_01172_),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08691_ (.I(_01173_),
    .Z(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08692_ (.I(_01174_),
    .Z(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08693_ (.I(_01175_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08694_ (.I(_01176_),
    .Z(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08695_ (.I(_01177_),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08696_ (.I0(\channels.exp_counter[0][0] ),
    .I1(\channels.exp_counter[1][0] ),
    .I2(\channels.exp_counter[2][0] ),
    .I3(\channels.exp_counter[3][0] ),
    .S0(_01162_),
    .S1(_01178_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08697_ (.I(_01175_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08698_ (.I(_01180_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08699_ (.I(_01181_),
    .Z(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08700_ (.I(_01182_),
    .Z(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08701_ (.I(_01183_),
    .Z(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08702_ (.I(_01162_),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08703_ (.I(_01185_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08704_ (.I0(\channels.exp_periods[0][0] ),
    .I1(\channels.exp_periods[1][0] ),
    .S(_01186_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08705_ (.I(_01185_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08706_ (.I(_01188_),
    .Z(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08707_ (.I(\channels.exp_periods[2][0] ),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08708_ (.A1(_01186_),
    .A2(\channels.exp_periods[3][0] ),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08709_ (.A1(_01189_),
    .A2(_01190_),
    .B(_01191_),
    .C(_01183_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08710_ (.A1(_01184_),
    .A2(_01187_),
    .B(_01192_),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08711_ (.A1(_01179_),
    .A2(_01193_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08712_ (.I0(\channels.exp_counter[0][2] ),
    .I1(\channels.exp_counter[1][2] ),
    .I2(\channels.exp_counter[2][2] ),
    .I3(\channels.exp_counter[3][2] ),
    .S0(_01185_),
    .S1(_01182_),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08713_ (.I(_01195_),
    .Z(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08714_ (.I(_01188_),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08715_ (.I(_01183_),
    .Z(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08716_ (.I0(\channels.exp_periods[0][2] ),
    .I1(\channels.exp_periods[1][2] ),
    .I2(\channels.exp_periods[2][2] ),
    .I3(\channels.exp_periods[3][2] ),
    .S0(_01197_),
    .S1(_01198_),
    .Z(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08717_ (.A1(_01196_),
    .A2(_01199_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08718_ (.I0(\channels.exp_counter[0][4] ),
    .I1(\channels.exp_counter[1][4] ),
    .I2(\channels.exp_counter[2][4] ),
    .I3(\channels.exp_counter[3][4] ),
    .S0(_01185_),
    .S1(_01182_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08719_ (.I0(\channels.exp_periods[0][4] ),
    .I1(\channels.exp_periods[1][4] ),
    .S(_01188_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08720_ (.I(\channels.exp_periods[2][4] ),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08721_ (.A1(_01186_),
    .A2(\channels.exp_periods[3][4] ),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08722_ (.A1(_01189_),
    .A2(_01203_),
    .B(_01204_),
    .C(_01183_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08723_ (.A1(_01184_),
    .A2(_01202_),
    .B(_01205_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08724_ (.A1(_01201_),
    .A2(_01206_),
    .Z(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08725_ (.I0(\channels.exp_counter[0][3] ),
    .I1(\channels.exp_counter[1][3] ),
    .I2(\channels.exp_counter[2][3] ),
    .I3(\channels.exp_counter[3][3] ),
    .S0(_01188_),
    .S1(_01182_),
    .Z(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08726_ (.I(_01208_),
    .Z(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08727_ (.I0(\channels.exp_periods[0][3] ),
    .I1(\channels.exp_periods[1][3] ),
    .S(_01197_),
    .Z(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08728_ (.I(_01186_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08729_ (.I(\channels.exp_periods[2][3] ),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08730_ (.A1(_01189_),
    .A2(\channels.exp_periods[3][3] ),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08731_ (.A1(_01211_),
    .A2(_01212_),
    .B(_01213_),
    .C(_01198_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08732_ (.A1(_01184_),
    .A2(_01210_),
    .B(_01214_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08733_ (.I0(\channels.exp_counter[0][1] ),
    .I1(\channels.exp_counter[1][1] ),
    .I2(\channels.exp_counter[2][1] ),
    .I3(\channels.exp_counter[3][1] ),
    .S0(_01162_),
    .S1(_01178_),
    .Z(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08734_ (.I0(\channels.exp_periods[0][1] ),
    .I1(\channels.exp_periods[1][1] ),
    .S(_01197_),
    .Z(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08735_ (.I(\channels.exp_periods[2][1] ),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08736_ (.A1(_01197_),
    .A2(\channels.exp_periods[3][1] ),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08737_ (.A1(_01189_),
    .A2(_01218_),
    .B(_01219_),
    .C(_01198_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08738_ (.A1(_01184_),
    .A2(_01217_),
    .B(_01220_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08739_ (.A1(_01209_),
    .A2(_01215_),
    .B1(_01216_),
    .B2(_01221_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08740_ (.A1(_01209_),
    .A2(_01215_),
    .B1(_01216_),
    .B2(_01221_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08741_ (.I(_01223_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08742_ (.A1(_01207_),
    .A2(_01222_),
    .A3(_01224_),
    .ZN(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08743_ (.A1(_01194_),
    .A2(_01200_),
    .A3(_01225_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08744_ (.I(_01226_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08745_ (.A1(_01179_),
    .A2(_01227_),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08746_ (.I(_01111_),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08747_ (.I(_01229_),
    .Z(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08748_ (.A1(\channels.exp_counter[1][0] ),
    .A2(_01115_),
    .B1(_01228_),
    .B2(_01230_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08749_ (.I(_01231_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08750_ (.A1(_01179_),
    .A2(_01216_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08751_ (.A1(_01179_),
    .A2(_01216_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08752_ (.A1(_01232_),
    .A2(_01233_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08753_ (.A1(_01227_),
    .A2(_01234_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08754_ (.A1(\channels.exp_counter[1][1] ),
    .A2(_01115_),
    .B1(_01235_),
    .B2(_01230_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08755_ (.I(_01236_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08756_ (.A1(_01196_),
    .A2(_01232_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08757_ (.A1(_01227_),
    .A2(_01237_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08758_ (.A1(\channels.exp_counter[1][2] ),
    .A2(_01115_),
    .B1(_01238_),
    .B2(_01230_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08759_ (.I(_01239_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08760_ (.I(_01113_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08761_ (.I(_01232_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08762_ (.A1(_01196_),
    .A2(_01209_),
    .A3(_01241_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08763_ (.A1(_01196_),
    .A2(_01241_),
    .B(_01209_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08764_ (.A1(_01226_),
    .A2(_01243_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08765_ (.A1(_01242_),
    .A2(_01244_),
    .Z(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08766_ (.A1(\channels.exp_counter[1][3] ),
    .A2(_01240_),
    .B1(_01245_),
    .B2(_01230_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08767_ (.I(_01246_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08768_ (.A1(_01201_),
    .A2(_01242_),
    .Z(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08769_ (.A1(_01227_),
    .A2(_01247_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08770_ (.A1(\channels.exp_counter[1][4] ),
    .A2(_01240_),
    .B1(_01248_),
    .B2(_01112_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08771_ (.I(_01249_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08772_ (.I(_01094_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08773_ (.I(_01250_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08774_ (.A1(\channels.exp_counter[2][0] ),
    .A2(_01101_),
    .B1(_01228_),
    .B2(_01251_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08775_ (.I(_01252_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08776_ (.A1(\channels.exp_counter[2][1] ),
    .A2(_01101_),
    .B1(_01235_),
    .B2(_01251_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08777_ (.I(_01253_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08778_ (.A1(\channels.exp_counter[2][2] ),
    .A2(_01101_),
    .B1(_01238_),
    .B2(_01251_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08779_ (.I(_01254_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08780_ (.I(_01099_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08781_ (.A1(\channels.exp_counter[2][3] ),
    .A2(_01255_),
    .B1(_01245_),
    .B2(_01251_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08782_ (.I(_01256_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08783_ (.A1(\channels.exp_counter[2][4] ),
    .A2(_01255_),
    .B1(_01248_),
    .B2(_01095_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08784_ (.I(_01257_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08785_ (.I(\channels.clk_div[2] ),
    .Z(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08786_ (.I(_01258_),
    .Z(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08787_ (.I(_01083_),
    .Z(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08788_ (.A1(_01259_),
    .A2(_01260_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08789_ (.I(_01261_),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08790_ (.A1(_01106_),
    .A2(_01262_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08791_ (.I(_01263_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08792_ (.I(_01264_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08793_ (.A1(_01098_),
    .A2(_01263_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08794_ (.I(_01266_),
    .Z(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08795_ (.I(_01267_),
    .Z(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08796_ (.A1(_01097_),
    .A2(_01265_),
    .B1(_01268_),
    .B2(\channels.ring_outs[0] ),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08797_ (.I(_01269_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08798_ (.I(\channels.accum[0][0] ),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08799_ (.I(_01266_),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08800_ (.I(_01271_),
    .Z(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08801_ (.I(_01260_),
    .Z(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08802_ (.I(_01273_),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08803_ (.I(_01107_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08804_ (.I(_01275_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08805_ (.I(_01276_),
    .Z(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08806_ (.A1(_01277_),
    .A2(\channels.ctrl_reg2[3] ),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08807_ (.A1(_01277_),
    .A2(\channels.ctrl_reg3[3] ),
    .B1(\channels.ctrl_reg1[3] ),
    .B2(_01262_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08808_ (.A1(_01274_),
    .A2(_01278_),
    .B(_01279_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08809_ (.A1(\channels.ctrl_reg3[1] ),
    .A2(\channels.sync_outs[1] ),
    .A3(_01093_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08810_ (.I(\channels.clk_div[1] ),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08811_ (.A1(_01258_),
    .A2(_01282_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08812_ (.I(_01283_),
    .Z(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08813_ (.I(_01284_),
    .Z(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08814_ (.I(_01285_),
    .Z(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08815_ (.I(_01286_),
    .Z(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08816_ (.I(_01287_),
    .Z(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08817_ (.I(_01288_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08818_ (.I(_01289_),
    .Z(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08819_ (.I(_01290_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08820_ (.I(_01291_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08821_ (.A1(\channels.ctrl_reg2[1] ),
    .A2(\channels.sync_outs[0] ),
    .A3(_01292_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08822_ (.A1(_01258_),
    .A2(\channels.clk_div[1] ),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08823_ (.I(_01294_),
    .Z(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08824_ (.I(_01295_),
    .Z(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08825_ (.I(_01296_),
    .Z(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08826_ (.I(_01297_),
    .Z(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08827_ (.I(_01298_),
    .Z(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08828_ (.I(_01299_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08829_ (.I(_01300_),
    .Z(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08830_ (.I(_01301_),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08831_ (.I(_01302_),
    .Z(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08832_ (.I(_01303_),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08833_ (.I(_01304_),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08834_ (.A1(\channels.ctrl_reg1[1] ),
    .A2(\channels.sync_outs[2] ),
    .A3(_01305_),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08835_ (.A1(_01281_),
    .A2(_01293_),
    .A3(_01306_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08836_ (.A1(_01280_),
    .A2(_01307_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08837_ (.I(_01308_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08838_ (.I(_01309_),
    .Z(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08839_ (.A1(\channels.freq3[0] ),
    .A2(_01085_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08840_ (.A1(\channels.freq2[0] ),
    .A2(_01284_),
    .B1(_01297_),
    .B2(\channels.freq1[0] ),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08841_ (.A1(_01311_),
    .A2(_01312_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08842_ (.I(_01198_),
    .Z(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08843_ (.I(_01152_),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08844_ (.I(_01315_),
    .Z(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08845_ (.I(_01316_),
    .Z(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08846_ (.I(_01317_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08847_ (.A1(_01318_),
    .A2(\channels.accum[1][0] ),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08848_ (.A1(_01156_),
    .A2(_01270_),
    .B(_01319_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08849_ (.I(\channels.accum[2][0] ),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08850_ (.A1(_01318_),
    .A2(\channels.accum[3][0] ),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08851_ (.A1(_01318_),
    .A2(_01321_),
    .B(_01322_),
    .C(_01169_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08852_ (.A1(_01314_),
    .A2(_01320_),
    .B(_01323_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08853_ (.A1(_01313_),
    .A2(_01324_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08854_ (.A1(_01310_),
    .A2(_01325_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08855_ (.I(_01263_),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08856_ (.I(_01327_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08857_ (.A1(_01270_),
    .A2(_01272_),
    .B1(_01326_),
    .B2(_01328_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08858_ (.I(_01305_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08859_ (.A1(_01081_),
    .A2(_01329_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08860_ (.I(_01330_),
    .Z(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08861_ (.I(_01331_),
    .Z(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08862_ (.I(_01308_),
    .Z(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08863_ (.A1(_01170_),
    .A2(_01320_),
    .B(_01323_),
    .C(_01313_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08864_ (.A1(\channels.freq3[1] ),
    .A2(_01085_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08865_ (.A1(\channels.freq2[1] ),
    .A2(_01284_),
    .B1(_01297_),
    .B2(\channels.freq1[1] ),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08866_ (.A1(_01335_),
    .A2(_01336_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08867_ (.I(_01168_),
    .Z(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08868_ (.I0(\channels.accum[0][1] ),
    .I1(\channels.accum[1][1] ),
    .I2(\channels.accum[2][1] ),
    .I3(\channels.accum[3][1] ),
    .S0(_01317_),
    .S1(_01338_),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08869_ (.A1(_01337_),
    .A2(_01339_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08870_ (.A1(_01334_),
    .A2(_01340_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08871_ (.A1(_01334_),
    .A2(_01340_),
    .Z(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08872_ (.A1(_01333_),
    .A2(_01341_),
    .A3(_01342_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08873_ (.I(_01266_),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08874_ (.A1(\channels.accum[0][1] ),
    .A2(_01344_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08875_ (.A1(_01332_),
    .A2(_01343_),
    .B(_01345_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08876_ (.I(\channels.accum[0][2] ),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08877_ (.I(_01309_),
    .Z(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08878_ (.A1(_01337_),
    .A2(_01339_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08879_ (.A1(\channels.freq3[2] ),
    .A2(_01086_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08880_ (.A1(\channels.freq2[2] ),
    .A2(_01285_),
    .B1(_01297_),
    .B2(\channels.freq1[2] ),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08881_ (.A1(_01349_),
    .A2(_01350_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08882_ (.I0(\channels.accum[0][2] ),
    .I1(\channels.accum[1][2] ),
    .I2(\channels.accum[2][2] ),
    .I3(\channels.accum[3][2] ),
    .S0(_01155_),
    .S1(_01169_),
    .Z(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08883_ (.A1(_01351_),
    .A2(_01352_),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08884_ (.A1(_01348_),
    .A2(_01342_),
    .A3(_01353_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08885_ (.A1(_01348_),
    .A2(_01342_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08886_ (.I(_01353_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08887_ (.A1(_01355_),
    .A2(_01356_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08888_ (.A1(_01347_),
    .A2(_01354_),
    .A3(_01357_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08889_ (.A1(_01346_),
    .A2(_01272_),
    .B1(_01358_),
    .B2(_01328_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08890_ (.I(_01309_),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08891_ (.A1(_01351_),
    .A2(_01352_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08892_ (.A1(_01360_),
    .A2(_01357_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08893_ (.A1(\channels.freq3[3] ),
    .A2(_01086_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08894_ (.A1(\channels.freq2[3] ),
    .A2(_01285_),
    .B1(_01298_),
    .B2(\channels.freq1[3] ),
    .ZN(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08895_ (.A1(_01362_),
    .A2(_01363_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08896_ (.I0(\channels.accum[0][3] ),
    .I1(\channels.accum[1][3] ),
    .I2(\channels.accum[2][3] ),
    .I3(\channels.accum[3][3] ),
    .S0(_01318_),
    .S1(_01170_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08897_ (.A1(_01364_),
    .A2(_01365_),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08898_ (.I(_01366_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08899_ (.A1(_01361_),
    .A2(_01367_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08900_ (.A1(_01359_),
    .A2(_01368_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08901_ (.I(_01267_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08902_ (.A1(\channels.accum[0][3] ),
    .A2(_01370_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08903_ (.A1(_01332_),
    .A2(_01369_),
    .B(_01371_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08904_ (.I(\channels.accum[0][4] ),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08905_ (.A1(_01360_),
    .A2(_01357_),
    .B(_01366_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08906_ (.A1(_01364_),
    .A2(_01365_),
    .B(_01373_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08907_ (.A1(\channels.freq3[4] ),
    .A2(_01086_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08908_ (.A1(\channels.freq2[4] ),
    .A2(_01285_),
    .B1(_01298_),
    .B2(\channels.freq1[4] ),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08909_ (.A1(_01375_),
    .A2(_01376_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08910_ (.I0(\channels.accum[0][4] ),
    .I1(\channels.accum[1][4] ),
    .I2(\channels.accum[2][4] ),
    .I3(\channels.accum[3][4] ),
    .S0(_01156_),
    .S1(_01171_),
    .Z(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08911_ (.A1(_01377_),
    .A2(_01378_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08912_ (.A1(_01374_),
    .A2(_01379_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08913_ (.A1(_01374_),
    .A2(_01379_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08914_ (.A1(_01347_),
    .A2(_01380_),
    .A3(_01381_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08915_ (.A1(_01372_),
    .A2(_01272_),
    .B1(_01382_),
    .B2(_01328_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08916_ (.A1(_01377_),
    .A2(_01378_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08917_ (.A1(_01383_),
    .A2(_01381_),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08918_ (.A1(\channels.freq3[5] ),
    .A2(_01087_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08919_ (.A1(\channels.freq2[5] ),
    .A2(_01286_),
    .B1(_01298_),
    .B2(\channels.freq1[5] ),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08920_ (.A1(_01385_),
    .A2(_01386_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08921_ (.I0(\channels.accum[0][5] ),
    .I1(\channels.accum[1][5] ),
    .I2(\channels.accum[2][5] ),
    .I3(\channels.accum[3][5] ),
    .S0(_01157_),
    .S1(_01171_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08922_ (.A1(_01387_),
    .A2(_01388_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08923_ (.A1(_01384_),
    .A2(_01389_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08924_ (.A1(_01359_),
    .A2(_01390_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08925_ (.A1(\channels.accum[0][5] ),
    .A2(_01370_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08926_ (.A1(_01332_),
    .A2(_01391_),
    .B(_01392_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08927_ (.I(\channels.accum[0][6] ),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08928_ (.A1(_01387_),
    .A2(_01388_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08929_ (.I(_01394_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08930_ (.A1(_01383_),
    .A2(_01381_),
    .B(_01389_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08931_ (.A1(\channels.freq3[6] ),
    .A2(_01087_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08932_ (.A1(\channels.freq2[6] ),
    .A2(_01286_),
    .B1(_01299_),
    .B2(\channels.freq1[6] ),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08933_ (.A1(_01397_),
    .A2(_01398_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08934_ (.I0(\channels.accum[0][6] ),
    .I1(\channels.accum[1][6] ),
    .I2(\channels.accum[2][6] ),
    .I3(\channels.accum[3][6] ),
    .S0(_01157_),
    .S1(_01172_),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08935_ (.A1(_01399_),
    .A2(_01400_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08936_ (.I(_01401_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08937_ (.A1(_01395_),
    .A2(_01396_),
    .A3(_01402_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08938_ (.A1(_01395_),
    .A2(_01396_),
    .B(_01402_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08939_ (.A1(_01347_),
    .A2(_01403_),
    .A3(_01404_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08940_ (.A1(_01393_),
    .A2(_01272_),
    .B1(_01405_),
    .B2(_01328_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08941_ (.A1(_01399_),
    .A2(_01400_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08942_ (.I(_01087_),
    .Z(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08943_ (.A1(\channels.freq3[7] ),
    .A2(_01407_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08944_ (.A1(\channels.freq2[7] ),
    .A2(_01287_),
    .B1(_01299_),
    .B2(\channels.freq1[7] ),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08945_ (.A1(_01408_),
    .A2(_01409_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08946_ (.I0(\channels.accum[0][7] ),
    .I1(\channels.accum[1][7] ),
    .I2(\channels.accum[2][7] ),
    .I3(\channels.accum[3][7] ),
    .S0(_01158_),
    .S1(_01173_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08947_ (.A1(_01410_),
    .A2(_01411_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08948_ (.A1(_01406_),
    .A2(_01404_),
    .A3(_01412_),
    .Z(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08949_ (.A1(_01406_),
    .A2(_01404_),
    .B(_01412_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08950_ (.A1(_01413_),
    .A2(_01414_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08951_ (.A1(_01359_),
    .A2(_01415_),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08952_ (.A1(\channels.accum[0][7] ),
    .A2(_01370_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08953_ (.A1(_01332_),
    .A2(_01416_),
    .B(_01417_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08954_ (.I(\channels.accum[0][8] ),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08955_ (.I(_01267_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08956_ (.A1(_01410_),
    .A2(_01411_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08957_ (.I(_01420_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08958_ (.A1(\channels.freq3[8] ),
    .A2(_01407_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08959_ (.A1(\channels.freq2[8] ),
    .A2(_01287_),
    .B1(_01299_),
    .B2(\channels.freq1[8] ),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08960_ (.A1(_01422_),
    .A2(_01423_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08961_ (.I0(\channels.accum[0][8] ),
    .I1(\channels.accum[1][8] ),
    .I2(\channels.accum[2][8] ),
    .I3(\channels.accum[3][8] ),
    .S0(_01158_),
    .S1(_01173_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08962_ (.A1(_01424_),
    .A2(_01425_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08963_ (.I(_01426_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08964_ (.A1(_01421_),
    .A2(_01414_),
    .A3(_01427_),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08965_ (.A1(_01421_),
    .A2(_01414_),
    .B(_01427_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08966_ (.A1(_01347_),
    .A2(_01428_),
    .A3(_01429_),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08967_ (.I(_01264_),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08968_ (.A1(_01418_),
    .A2(_01419_),
    .B1(_01430_),
    .B2(_01431_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08969_ (.I(_01331_),
    .Z(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08970_ (.A1(_01424_),
    .A2(_01425_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08971_ (.A1(\channels.freq3[9] ),
    .A2(_01088_),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08972_ (.I(_01286_),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08973_ (.A1(\channels.freq2[9] ),
    .A2(_01435_),
    .B1(_01300_),
    .B2(\channels.freq1[9] ),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08974_ (.A1(_01434_),
    .A2(_01436_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _08975_ (.I0(\channels.accum[0][9] ),
    .I1(\channels.accum[1][9] ),
    .I2(\channels.accum[2][9] ),
    .I3(\channels.accum[3][9] ),
    .S0(_01158_),
    .S1(_01173_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08976_ (.A1(_01437_),
    .A2(_01438_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08977_ (.A1(_01433_),
    .A2(_01429_),
    .A3(_01439_),
    .Z(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08978_ (.A1(_01433_),
    .A2(_01429_),
    .B(_01439_),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08979_ (.A1(_01440_),
    .A2(_01441_),
    .ZN(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08980_ (.A1(_01359_),
    .A2(_01442_),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08981_ (.A1(\channels.accum[0][9] ),
    .A2(_01370_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08982_ (.A1(_01432_),
    .A2(_01443_),
    .B(_01444_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08983_ (.I(\channels.accum[0][10] ),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08984_ (.I(_01308_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08985_ (.A1(_01437_),
    .A2(_01438_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08986_ (.I(_01447_),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08987_ (.I(_01407_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08988_ (.A1(\channels.freq3[10] ),
    .A2(_01449_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08989_ (.A1(\channels.freq2[10] ),
    .A2(_01288_),
    .B1(_01300_),
    .B2(\channels.freq1[10] ),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08990_ (.A1(_01450_),
    .A2(_01451_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08991_ (.I0(\channels.accum[0][10] ),
    .I1(\channels.accum[1][10] ),
    .I2(\channels.accum[2][10] ),
    .I3(\channels.accum[3][10] ),
    .S0(_01159_),
    .S1(_01174_),
    .Z(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08992_ (.A1(_01452_),
    .A2(_01453_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08993_ (.I(_01454_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08994_ (.A1(_01448_),
    .A2(_01441_),
    .A3(_01455_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08995_ (.A1(_01448_),
    .A2(_01441_),
    .B(_01455_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08996_ (.A1(_01446_),
    .A2(_01456_),
    .A3(_01457_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08997_ (.A1(_01445_),
    .A2(_01419_),
    .B1(_01458_),
    .B2(_01431_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08998_ (.I(_01309_),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08999_ (.A1(_01452_),
    .A2(_01453_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09000_ (.A1(\channels.freq3[11] ),
    .A2(_01090_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09001_ (.A1(\channels.freq2[11] ),
    .A2(_01289_),
    .B1(_01302_),
    .B2(\channels.freq1[11] ),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09002_ (.A1(_01461_),
    .A2(_01462_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _09003_ (.I0(\channels.accum[0][11] ),
    .I1(\channels.accum[1][11] ),
    .I2(\channels.accum[2][11] ),
    .I3(\channels.accum[3][11] ),
    .S0(_01159_),
    .S1(_01175_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09004_ (.A1(_01463_),
    .A2(_01464_),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09005_ (.A1(_01460_),
    .A2(_01457_),
    .A3(_01465_),
    .Z(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09006_ (.A1(_01460_),
    .A2(_01457_),
    .B(_01465_),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09007_ (.A1(_01466_),
    .A2(_01467_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09008_ (.A1(_01459_),
    .A2(_01468_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09009_ (.I(_01266_),
    .Z(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09010_ (.I(_01470_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09011_ (.A1(\channels.accum[0][11] ),
    .A2(_01471_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09012_ (.A1(_01432_),
    .A2(_01469_),
    .B(_01472_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09013_ (.I(\channels.accum[0][12] ),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09014_ (.A1(_01463_),
    .A2(_01464_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09015_ (.I(_01474_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09016_ (.A1(\channels.freq3[12] ),
    .A2(_01090_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09017_ (.A1(\channels.freq2[12] ),
    .A2(_01289_),
    .B1(_01302_),
    .B2(\channels.freq1[12] ),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09018_ (.A1(_01476_),
    .A2(_01477_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09019_ (.I0(\channels.accum[0][12] ),
    .I1(\channels.accum[1][12] ),
    .I2(\channels.accum[2][12] ),
    .I3(\channels.accum[3][12] ),
    .S0(_01150_),
    .S1(_01164_),
    .Z(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09020_ (.I(_01479_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09021_ (.A1(_01478_),
    .A2(_01480_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09022_ (.I(_01481_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09023_ (.A1(_01475_),
    .A2(_01467_),
    .A3(_01482_),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09024_ (.A1(_01475_),
    .A2(_01467_),
    .B(_01482_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09025_ (.A1(_01446_),
    .A2(_01483_),
    .A3(_01484_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09026_ (.A1(_01473_),
    .A2(_01419_),
    .B1(_01485_),
    .B2(_01431_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09027_ (.A1(_01478_),
    .A2(_01480_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09028_ (.A1(\channels.freq3[13] ),
    .A2(_01090_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09029_ (.A1(\channels.freq2[13] ),
    .A2(_01289_),
    .B1(_01303_),
    .B2(\channels.freq1[13] ),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09030_ (.A1(_01487_),
    .A2(_01488_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09031_ (.I(_00010_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09032_ (.I0(\channels.accum[0][13] ),
    .I1(\channels.accum[1][13] ),
    .I2(\channels.accum[2][13] ),
    .I3(\channels.accum[3][13] ),
    .S0(_01148_),
    .S1(_01490_),
    .Z(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09033_ (.I(_01491_),
    .Z(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09034_ (.A1(_01489_),
    .A2(_01492_),
    .ZN(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09035_ (.A1(_01486_),
    .A2(_01484_),
    .A3(_01493_),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09036_ (.A1(_01486_),
    .A2(_01484_),
    .B(_01493_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09037_ (.A1(_01494_),
    .A2(_01495_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09038_ (.A1(_01459_),
    .A2(_01496_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09039_ (.A1(\channels.accum[0][13] ),
    .A2(_01471_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09040_ (.A1(_01432_),
    .A2(_01497_),
    .B(_01498_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09041_ (.I(\channels.accum[0][14] ),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09042_ (.A1(_01489_),
    .A2(_01492_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09043_ (.I(_01500_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09044_ (.A1(\channels.freq3[14] ),
    .A2(_01091_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09045_ (.A1(\channels.freq2[14] ),
    .A2(_01290_),
    .B1(_01303_),
    .B2(\channels.freq1[14] ),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09046_ (.A1(_01502_),
    .A2(_01503_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09047_ (.I(_01148_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09048_ (.I(_01163_),
    .Z(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09049_ (.I0(\channels.accum[0][14] ),
    .I1(\channels.accum[1][14] ),
    .I2(\channels.accum[2][14] ),
    .I3(\channels.accum[3][14] ),
    .S0(_01505_),
    .S1(_01506_),
    .Z(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09050_ (.I(_01507_),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09051_ (.A1(_01504_),
    .A2(_01508_),
    .Z(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09052_ (.I(_01509_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09053_ (.A1(_01501_),
    .A2(_01495_),
    .A3(_01510_),
    .Z(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09054_ (.A1(_01501_),
    .A2(_01495_),
    .B(_01510_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09055_ (.A1(_01446_),
    .A2(_01511_),
    .A3(_01512_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09056_ (.A1(_01499_),
    .A2(_01419_),
    .B1(_01513_),
    .B2(_01431_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09057_ (.A1(_01504_),
    .A2(_01507_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09058_ (.A1(\channels.freq3[15] ),
    .A2(_01091_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09059_ (.A1(\channels.freq2[15] ),
    .A2(_01290_),
    .B1(_01303_),
    .B2(\channels.freq1[15] ),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09060_ (.A1(_01515_),
    .A2(_01516_),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09061_ (.I0(\channels.accum[0][15] ),
    .I1(\channels.accum[1][15] ),
    .I2(\channels.accum[2][15] ),
    .I3(\channels.accum[3][15] ),
    .S0(_00009_),
    .S1(_01163_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09062_ (.I(_01518_),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09063_ (.I(_01519_),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09064_ (.A1(_01517_),
    .A2(_01520_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09065_ (.A1(_01514_),
    .A2(_01512_),
    .A3(_01521_),
    .Z(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09066_ (.A1(_01514_),
    .A2(_01512_),
    .B(_01521_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09067_ (.A1(_01522_),
    .A2(_01523_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09068_ (.A1(_01459_),
    .A2(_01524_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09069_ (.A1(\channels.accum[0][15] ),
    .A2(_01471_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09070_ (.A1(_01432_),
    .A2(_01525_),
    .B(_01526_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09071_ (.I(\channels.accum[0][16] ),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09072_ (.I(_01267_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09073_ (.A1(_01515_),
    .A2(_01516_),
    .B(_01520_),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09074_ (.I0(\channels.accum[0][16] ),
    .I1(\channels.accum[1][16] ),
    .I2(\channels.accum[2][16] ),
    .I3(\channels.accum[3][16] ),
    .S0(_01149_),
    .S1(_01490_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09075_ (.I(_01530_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09076_ (.A1(_01529_),
    .A2(_01523_),
    .A3(_01531_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09077_ (.A1(_01529_),
    .A2(_01523_),
    .B(_01531_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09078_ (.A1(_01446_),
    .A2(_01532_),
    .A3(_01533_),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09079_ (.I(_01264_),
    .Z(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09080_ (.A1(_01527_),
    .A2(_01528_),
    .B1(_01534_),
    .B2(_01535_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09081_ (.I(_01533_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09082_ (.I0(\channels.accum[0][17] ),
    .I1(\channels.accum[1][17] ),
    .I2(\channels.accum[2][17] ),
    .I3(\channels.accum[3][17] ),
    .S0(_01149_),
    .S1(_01490_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09083_ (.I(_01537_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09084_ (.A1(_01536_),
    .A2(_01538_),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09085_ (.A1(_01333_),
    .A2(_01539_),
    .Z(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09086_ (.A1(\channels.accum[0][17] ),
    .A2(_01344_),
    .B1(_01540_),
    .B2(_01265_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09087_ (.I(_01541_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09088_ (.I(\channels.accum[0][18] ),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09089_ (.I0(\channels.accum[0][18] ),
    .I1(\channels.accum[1][18] ),
    .I2(\channels.accum[2][18] ),
    .I3(\channels.accum[3][18] ),
    .S0(_01505_),
    .S1(_01506_),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09090_ (.I(_01543_),
    .Z(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09091_ (.A1(_01536_),
    .A2(_01538_),
    .B(_01544_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09092_ (.A1(_01536_),
    .A2(_01538_),
    .A3(_01544_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09093_ (.I(_01546_),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09094_ (.A1(_01333_),
    .A2(_01547_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09095_ (.A1(_01545_),
    .A2(_01548_),
    .Z(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09096_ (.A1(_01542_),
    .A2(_01528_),
    .B1(_01549_),
    .B2(_01535_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09097_ (.I(_01331_),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09098_ (.I0(\channels.accum[0][19] ),
    .I1(\channels.accum[1][19] ),
    .I2(\channels.accum[2][19] ),
    .I3(\channels.accum[3][19] ),
    .S0(_01505_),
    .S1(_01506_),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09099_ (.I(_01551_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09100_ (.I(_01552_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09101_ (.A1(_01547_),
    .A2(_01553_),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09102_ (.A1(_01459_),
    .A2(_01554_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09103_ (.A1(\channels.accum[0][19] ),
    .A2(_01471_),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09104_ (.A1(_01550_),
    .A2(_01555_),
    .B(_01556_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09105_ (.I(\channels.accum[0][20] ),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09106_ (.A1(_01547_),
    .A2(_01553_),
    .ZN(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09107_ (.I0(\channels.accum[0][20] ),
    .I1(\channels.accum[1][20] ),
    .I2(\channels.accum[2][20] ),
    .I3(\channels.accum[3][20] ),
    .S0(_01148_),
    .S1(_01163_),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09108_ (.I(_01559_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09109_ (.A1(_01558_),
    .A2(_01560_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09110_ (.A1(_01310_),
    .A2(_01561_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09111_ (.A1(_01557_),
    .A2(_01528_),
    .B1(_01562_),
    .B2(_01535_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09112_ (.I(_01559_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09113_ (.A1(_01546_),
    .A2(_01553_),
    .A3(_01563_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09114_ (.I0(\channels.accum[0][21] ),
    .I1(\channels.accum[1][21] ),
    .I2(\channels.accum[2][21] ),
    .I3(\channels.accum[3][21] ),
    .S0(_01149_),
    .S1(_01490_),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09115_ (.I(_01565_),
    .Z(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09116_ (.A1(_01564_),
    .A2(_01566_),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09117_ (.A1(_01564_),
    .A2(_01566_),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09118_ (.A1(_01333_),
    .A2(_01567_),
    .A3(_01568_),
    .ZN(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09119_ (.I(_01470_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09120_ (.A1(\channels.accum[0][21] ),
    .A2(_01570_),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09121_ (.A1(_01550_),
    .A2(_01569_),
    .B(_01571_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09122_ (.I(\channels.accum[0][22] ),
    .ZN(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09123_ (.I(\channels.accum[1][22] ),
    .ZN(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09124_ (.I(\channels.accum[2][22] ),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09125_ (.I(\channels.accum[3][22] ),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09126_ (.I0(_01572_),
    .I1(_01573_),
    .I2(_01574_),
    .I3(_01575_),
    .S0(_01150_),
    .S1(_01164_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09127_ (.A1(_01568_),
    .A2(_01576_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09128_ (.A1(_01310_),
    .A2(_01577_),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09129_ (.A1(_01572_),
    .A2(_01528_),
    .B1(_01578_),
    .B2(_01535_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09130_ (.A1(_01568_),
    .A2(_01576_),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09131_ (.A1(_01097_),
    .A2(_01579_),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09132_ (.A1(_01310_),
    .A2(_01580_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09133_ (.A1(\channels.accum[0][23] ),
    .A2(_01570_),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09134_ (.A1(_01550_),
    .A2(_01581_),
    .B(_01582_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09135_ (.I(\channels.lfsr[0][17] ),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09136_ (.I(\channels.lfsr[1][17] ),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09137_ (.I(\channels.lfsr[2][17] ),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09138_ (.I(\channels.lfsr[3][17] ),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09139_ (.I0(_01583_),
    .I1(_01584_),
    .I2(_01585_),
    .I3(_01586_),
    .S0(_01211_),
    .S1(_01314_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _09140_ (.I0(\channels.lfsr[0][22] ),
    .I1(\channels.lfsr[1][22] ),
    .I2(\channels.lfsr[2][22] ),
    .I3(\channels.lfsr[3][22] ),
    .S0(_01211_),
    .S1(_01314_),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09141_ (.A1(_01587_),
    .A2(_01588_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09142_ (.A1(_01280_),
    .A2(_01589_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09143_ (.I(_01093_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09144_ (.I(_01259_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09145_ (.I(_01592_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09146_ (.A1(_01593_),
    .A2(_01274_),
    .B(_01106_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09147_ (.I(_01594_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09148_ (.I(_01595_),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09149_ (.A1(_01280_),
    .A2(_01547_),
    .A3(_01552_),
    .A4(_01596_),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09150_ (.A1(_01591_),
    .A2(_01597_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09151_ (.I(_01598_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09152_ (.I(_01040_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09153_ (.A1(_01600_),
    .A2(_01598_),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09154_ (.I(_01601_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09155_ (.I(_01602_),
    .Z(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09156_ (.I(\channels.lfsr[2][0] ),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09157_ (.A1(_01590_),
    .A2(_01599_),
    .B1(_01603_),
    .B2(_01604_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09158_ (.I(\channels.lfsr[2][1] ),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09159_ (.I(\channels.lfsr[0][0] ),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09160_ (.I(\channels.lfsr[1][0] ),
    .ZN(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09161_ (.I(\channels.lfsr[3][0] ),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09162_ (.I0(_01606_),
    .I1(_01607_),
    .I2(_01604_),
    .I3(_01608_),
    .S0(_01150_),
    .S1(_01164_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09163_ (.I(_01599_),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09164_ (.A1(_01605_),
    .A2(_01603_),
    .B1(_01609_),
    .B2(_01610_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09165_ (.I(\channels.lfsr[2][2] ),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09166_ (.I(\channels.lfsr[0][1] ),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09167_ (.I(\channels.lfsr[1][1] ),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09168_ (.I(\channels.lfsr[3][1] ),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09169_ (.I(_01211_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09170_ (.I(_01615_),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09171_ (.I(_01314_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09172_ (.I(_01617_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _09173_ (.I0(_01612_),
    .I1(_01613_),
    .I2(_01605_),
    .I3(_01614_),
    .S0(_01616_),
    .S1(_01618_),
    .Z(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09174_ (.A1(_01611_),
    .A2(_01603_),
    .B1(_01619_),
    .B2(_01610_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09175_ (.I(\channels.lfsr[2][3] ),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09176_ (.I(_01601_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09177_ (.I(_01621_),
    .Z(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09178_ (.I(\channels.lfsr[0][2] ),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09179_ (.I(\channels.lfsr[1][2] ),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09180_ (.I(\channels.lfsr[3][2] ),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09181_ (.I0(_01623_),
    .I1(_01624_),
    .I2(_01611_),
    .I3(_01625_),
    .S0(_01151_),
    .S1(_01165_),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09182_ (.A1(_01620_),
    .A2(_01622_),
    .B1(_01626_),
    .B2(_01610_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09183_ (.I(\channels.lfsr[2][4] ),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09184_ (.I(\channels.lfsr[0][3] ),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09185_ (.I(\channels.lfsr[1][3] ),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09186_ (.I(\channels.lfsr[3][3] ),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09187_ (.I0(_01628_),
    .I1(_01629_),
    .I2(_01620_),
    .I3(_01630_),
    .S0(_01616_),
    .S1(_01618_),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09188_ (.A1(_01627_),
    .A2(_01622_),
    .B1(_01631_),
    .B2(_01610_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09189_ (.I(\channels.lfsr[2][5] ),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09190_ (.I(\channels.lfsr[0][4] ),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09191_ (.I(\channels.lfsr[1][4] ),
    .ZN(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09192_ (.I(\channels.lfsr[3][4] ),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09193_ (.I0(_01633_),
    .I1(_01634_),
    .I2(_01627_),
    .I3(_01635_),
    .S0(_01616_),
    .S1(_01618_),
    .Z(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09194_ (.I(_01598_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09195_ (.I(_01637_),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09196_ (.A1(_01632_),
    .A2(_01622_),
    .B1(_01636_),
    .B2(_01638_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09197_ (.I(\channels.lfsr[2][6] ),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09198_ (.I(\channels.lfsr[0][5] ),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09199_ (.I(\channels.lfsr[1][5] ),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09200_ (.I(\channels.lfsr[3][5] ),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09201_ (.I0(_01640_),
    .I1(_01641_),
    .I2(_01632_),
    .I3(_01642_),
    .S0(_01151_),
    .S1(_01165_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09202_ (.A1(_01639_),
    .A2(_01622_),
    .B1(_01643_),
    .B2(_01638_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09203_ (.I(\channels.lfsr[2][7] ),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09204_ (.I(_01621_),
    .Z(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09205_ (.I(\channels.lfsr[0][6] ),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09206_ (.I(\channels.lfsr[1][6] ),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09207_ (.I(\channels.lfsr[3][6] ),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09208_ (.I0(_01646_),
    .I1(_01647_),
    .I2(_01639_),
    .I3(_01648_),
    .S0(_01616_),
    .S1(_01618_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09209_ (.A1(_01644_),
    .A2(_01645_),
    .B1(_01649_),
    .B2(_01638_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09210_ (.I(\channels.lfsr[2][8] ),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09211_ (.I(\channels.lfsr[0][7] ),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09212_ (.I(\channels.lfsr[1][7] ),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09213_ (.I(\channels.lfsr[3][7] ),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09214_ (.I(_01615_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09215_ (.I(_01617_),
    .Z(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09216_ (.I0(_01651_),
    .I1(_01652_),
    .I2(_01644_),
    .I3(_01653_),
    .S0(_01654_),
    .S1(_01655_),
    .Z(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09217_ (.A1(_01650_),
    .A2(_01645_),
    .B1(_01656_),
    .B2(_01638_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09218_ (.I(\channels.lfsr[2][9] ),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09219_ (.I(\channels.lfsr[0][8] ),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09220_ (.I(\channels.lfsr[1][8] ),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09221_ (.I(\channels.lfsr[3][8] ),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09222_ (.I0(_01658_),
    .I1(_01659_),
    .I2(_01650_),
    .I3(_01660_),
    .S0(_01654_),
    .S1(_01655_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09223_ (.I(_01637_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09224_ (.A1(_01657_),
    .A2(_01645_),
    .B1(_01661_),
    .B2(_01662_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09225_ (.I(\channels.lfsr[2][10] ),
    .ZN(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09226_ (.I(\channels.lfsr[0][9] ),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09227_ (.I(\channels.lfsr[1][9] ),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09228_ (.I(\channels.lfsr[3][9] ),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09229_ (.I(_01165_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09230_ (.I0(_01664_),
    .I1(_01665_),
    .I2(_01657_),
    .I3(_01666_),
    .S0(_01152_),
    .S1(_01667_),
    .Z(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09231_ (.A1(_01663_),
    .A2(_01645_),
    .B1(_01668_),
    .B2(_01662_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09232_ (.I(\channels.lfsr[2][11] ),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09233_ (.I(_01621_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09234_ (.I(\channels.lfsr[0][10] ),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09235_ (.I(\channels.lfsr[1][10] ),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09236_ (.I(\channels.lfsr[3][10] ),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09237_ (.I0(_01671_),
    .I1(_01672_),
    .I2(_01663_),
    .I3(_01673_),
    .S0(_01654_),
    .S1(_01655_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09238_ (.A1(_01669_),
    .A2(_01670_),
    .B1(_01674_),
    .B2(_01662_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09239_ (.I(\channels.lfsr[2][12] ),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09240_ (.I(\channels.lfsr[0][11] ),
    .ZN(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09241_ (.I(\channels.lfsr[1][11] ),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09242_ (.I(\channels.lfsr[3][11] ),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09243_ (.I0(_01676_),
    .I1(_01677_),
    .I2(_01669_),
    .I3(_01678_),
    .S0(_01315_),
    .S1(_01667_),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09244_ (.A1(_01675_),
    .A2(_01670_),
    .B1(_01679_),
    .B2(_01662_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09245_ (.I(\channels.lfsr[2][13] ),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09246_ (.I(\channels.lfsr[0][12] ),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09247_ (.I(\channels.lfsr[1][12] ),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09248_ (.I(\channels.lfsr[3][12] ),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09249_ (.I0(_01681_),
    .I1(_01682_),
    .I2(_01675_),
    .I3(_01683_),
    .S0(_01654_),
    .S1(_01655_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09250_ (.I(_01637_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09251_ (.A1(_01680_),
    .A2(_01670_),
    .B1(_01684_),
    .B2(_01685_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09252_ (.I(\channels.lfsr[2][14] ),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09253_ (.I(\channels.lfsr[0][13] ),
    .ZN(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09254_ (.I(\channels.lfsr[1][13] ),
    .ZN(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09255_ (.I(\channels.lfsr[3][13] ),
    .ZN(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09256_ (.I(_01615_),
    .Z(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09257_ (.I(_01617_),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09258_ (.I0(_01687_),
    .I1(_01688_),
    .I2(_01680_),
    .I3(_01689_),
    .S0(_01690_),
    .S1(_01691_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09259_ (.A1(_01686_),
    .A2(_01670_),
    .B1(_01692_),
    .B2(_01685_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09260_ (.I(\channels.lfsr[2][15] ),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09261_ (.I(_01621_),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09262_ (.I(\channels.lfsr[0][14] ),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09263_ (.I(\channels.lfsr[1][14] ),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09264_ (.I(\channels.lfsr[3][14] ),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09265_ (.I(_01667_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09266_ (.I(_01698_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09267_ (.I0(_01695_),
    .I1(_01696_),
    .I2(_01686_),
    .I3(_01697_),
    .S0(_01154_),
    .S1(_01699_),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09268_ (.A1(_01693_),
    .A2(_01694_),
    .B1(_01700_),
    .B2(_01685_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09269_ (.I(\channels.lfsr[2][16] ),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09270_ (.I(\channels.lfsr[0][15] ),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09271_ (.I(\channels.lfsr[1][15] ),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09272_ (.I(\channels.lfsr[3][15] ),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09273_ (.I0(_01702_),
    .I1(_01703_),
    .I2(_01693_),
    .I3(_01704_),
    .S0(_01690_),
    .S1(_01691_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09274_ (.A1(_01701_),
    .A2(_01694_),
    .B1(_01705_),
    .B2(_01685_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09275_ (.I(\channels.lfsr[0][16] ),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09276_ (.I(\channels.lfsr[1][16] ),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09277_ (.I(\channels.lfsr[3][16] ),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09278_ (.I0(_01706_),
    .I1(_01707_),
    .I2(_01701_),
    .I3(_01708_),
    .S0(_01690_),
    .S1(_01691_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09279_ (.I(_01637_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09280_ (.A1(_01585_),
    .A2(_01694_),
    .B1(_01709_),
    .B2(_01710_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09281_ (.I(\channels.lfsr[2][18] ),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09282_ (.A1(_01587_),
    .A2(_01599_),
    .B1(_01603_),
    .B2(_01711_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09283_ (.I(\channels.lfsr[2][19] ),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09284_ (.I(\channels.lfsr[0][18] ),
    .ZN(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09285_ (.I(\channels.lfsr[1][18] ),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09286_ (.I(\channels.lfsr[3][18] ),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09287_ (.I0(_01713_),
    .I1(_01714_),
    .I2(_01711_),
    .I3(_01715_),
    .S0(_01154_),
    .S1(_01168_),
    .Z(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09288_ (.A1(_01712_),
    .A2(_01694_),
    .B1(_01716_),
    .B2(_01710_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09289_ (.I(\channels.lfsr[2][20] ),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09290_ (.I(\channels.lfsr[0][19] ),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09291_ (.I(\channels.lfsr[1][19] ),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09292_ (.I(\channels.lfsr[3][19] ),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09293_ (.I0(_01718_),
    .I1(_01719_),
    .I2(_01712_),
    .I3(_01720_),
    .S0(_01690_),
    .S1(_01691_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09294_ (.A1(_01717_),
    .A2(_01602_),
    .B1(_01721_),
    .B2(_01710_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09295_ (.I(\channels.lfsr[2][21] ),
    .ZN(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09296_ (.I(\channels.lfsr[0][20] ),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09297_ (.I(\channels.lfsr[1][20] ),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09298_ (.I(\channels.lfsr[3][20] ),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09299_ (.I0(_01723_),
    .I1(_01724_),
    .I2(_01717_),
    .I3(_01725_),
    .S0(_01155_),
    .S1(_01338_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09300_ (.A1(_01722_),
    .A2(_01602_),
    .B1(_01726_),
    .B2(_01710_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09301_ (.I(\channels.lfsr[2][22] ),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09302_ (.I(\channels.lfsr[0][21] ),
    .ZN(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09303_ (.I(\channels.lfsr[1][21] ),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09304_ (.I(\channels.lfsr[3][21] ),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _09305_ (.I0(_01728_),
    .I1(_01729_),
    .I2(_01722_),
    .I3(_01730_),
    .S0(_01615_),
    .S1(_01617_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09306_ (.A1(_01727_),
    .A2(_01602_),
    .B1(_01731_),
    .B2(_01599_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09307_ (.A1(_01292_),
    .A2(_01597_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09308_ (.I(_01732_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09309_ (.I(_01733_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09310_ (.A1(_01600_),
    .A2(_01732_),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09311_ (.I(_01735_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09312_ (.I(_01736_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09313_ (.A1(_01590_),
    .A2(_01734_),
    .B1(_01737_),
    .B2(_01607_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09314_ (.A1(_01609_),
    .A2(_01734_),
    .B1(_01737_),
    .B2(_01613_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09315_ (.A1(_01619_),
    .A2(_01734_),
    .B1(_01737_),
    .B2(_01624_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09316_ (.A1(_01626_),
    .A2(_01734_),
    .B1(_01737_),
    .B2(_01629_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09317_ (.I(_01732_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09318_ (.I(_01738_),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09319_ (.I(_01735_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09320_ (.I(_01740_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09321_ (.A1(_01631_),
    .A2(_01739_),
    .B1(_01741_),
    .B2(_01634_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09322_ (.A1(_01636_),
    .A2(_01739_),
    .B1(_01741_),
    .B2(_01641_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09323_ (.A1(_01643_),
    .A2(_01739_),
    .B1(_01741_),
    .B2(_01647_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09324_ (.A1(_01649_),
    .A2(_01739_),
    .B1(_01741_),
    .B2(_01652_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09325_ (.I(_01738_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09326_ (.I(_01740_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09327_ (.A1(_01656_),
    .A2(_01742_),
    .B1(_01743_),
    .B2(_01659_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09328_ (.A1(_01661_),
    .A2(_01742_),
    .B1(_01743_),
    .B2(_01665_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09329_ (.A1(_01668_),
    .A2(_01742_),
    .B1(_01743_),
    .B2(_01672_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09330_ (.A1(_01674_),
    .A2(_01742_),
    .B1(_01743_),
    .B2(_01677_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09331_ (.I(_01738_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09332_ (.I(_01740_),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09333_ (.A1(_01679_),
    .A2(_01744_),
    .B1(_01745_),
    .B2(_01682_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09334_ (.A1(_01684_),
    .A2(_01744_),
    .B1(_01745_),
    .B2(_01688_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09335_ (.A1(_01692_),
    .A2(_01744_),
    .B1(_01745_),
    .B2(_01696_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09336_ (.A1(_01700_),
    .A2(_01744_),
    .B1(_01745_),
    .B2(_01703_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09337_ (.I(_01738_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09338_ (.I(_01740_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09339_ (.A1(_01705_),
    .A2(_01746_),
    .B1(_01747_),
    .B2(_01707_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09340_ (.A1(_01709_),
    .A2(_01746_),
    .B1(_01747_),
    .B2(_01584_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09341_ (.A1(_01587_),
    .A2(_01746_),
    .B1(_01747_),
    .B2(_01714_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09342_ (.A1(_01716_),
    .A2(_01746_),
    .B1(_01747_),
    .B2(_01719_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09343_ (.A1(_01721_),
    .A2(_01733_),
    .B1(_01736_),
    .B2(_01724_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09344_ (.A1(_01726_),
    .A2(_01733_),
    .B1(_01736_),
    .B2(_01729_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09345_ (.I(\channels.lfsr[1][22] ),
    .ZN(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09346_ (.A1(_01731_),
    .A2(_01733_),
    .B1(_01736_),
    .B2(_01748_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09347_ (.I(net7),
    .ZN(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09348_ (.I(_01749_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09349_ (.I(_01750_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09350_ (.I(_01751_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09351_ (.I(_01020_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09352_ (.I(\filters.filt_1 ),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09353_ (.I(_01754_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09354_ (.I(_01755_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09355_ (.I(_01756_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09356_ (.I(_01757_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09357_ (.I(_01020_),
    .Z(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09358_ (.I(_01071_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09359_ (.I(_01760_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09360_ (.I(_01761_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09361_ (.I(_01762_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09362_ (.A1(_01758_),
    .A2(_01759_),
    .B(_01763_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09363_ (.A1(_01752_),
    .A2(_01753_),
    .B(_01764_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09364_ (.I(net8),
    .ZN(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09365_ (.I(_01765_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09366_ (.I(_01766_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09367_ (.I(\filters.filt_2 ),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09368_ (.I(_01768_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09369_ (.I(_01769_),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09370_ (.I(_01770_),
    .Z(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09371_ (.I(_01771_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09372_ (.I(_01762_),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09373_ (.A1(_01772_),
    .A2(_01759_),
    .B(_01773_),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09374_ (.A1(_01767_),
    .A2(_01753_),
    .B(_01774_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09375_ (.I(net9),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09376_ (.I(_01775_),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09377_ (.I(_01776_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09378_ (.I(\filters.filt_3 ),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09379_ (.I(_01778_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09380_ (.I(_01779_),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09381_ (.I(_01780_),
    .Z(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09382_ (.I(_01781_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09383_ (.I(_01782_),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09384_ (.A1(_01783_),
    .A2(_01759_),
    .B(_01773_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09385_ (.A1(_01777_),
    .A2(_01753_),
    .B(_01784_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09386_ (.I(net10),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09387_ (.I(_01785_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09388_ (.I(_01786_),
    .Z(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09389_ (.A1(\filters.res_filt[3] ),
    .A2(_01759_),
    .B(_01773_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09390_ (.A1(_01787_),
    .A2(_01753_),
    .B(_01788_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09391_ (.I(_01016_),
    .Z(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09392_ (.I(_01789_),
    .Z(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09393_ (.I(_01790_),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09394_ (.I(_01011_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09395_ (.A1(net2),
    .A2(net1),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09396_ (.A1(_01792_),
    .A2(_01793_),
    .Z(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09397_ (.A1(_01012_),
    .A2(net3),
    .A3(_01794_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09398_ (.I(_01795_),
    .Z(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09399_ (.A1(_01791_),
    .A2(_01796_),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09400_ (.I(_01797_),
    .Z(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09401_ (.I(_01797_),
    .Z(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09402_ (.A1(\filters.mode_vol[0] ),
    .A2(_01799_),
    .B(_01773_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09403_ (.A1(_01752_),
    .A2(_01798_),
    .B(_01800_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09404_ (.I(_01762_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09405_ (.A1(\filters.mode_vol[1] ),
    .A2(_01799_),
    .B(_01801_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09406_ (.A1(_01767_),
    .A2(_01798_),
    .B(_01802_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09407_ (.A1(\filters.mode_vol[2] ),
    .A2(_01799_),
    .B(_01801_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09408_ (.A1(_01777_),
    .A2(_01798_),
    .B(_01803_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09409_ (.A1(\filters.mode_vol[3] ),
    .A2(_01799_),
    .B(_01801_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09410_ (.A1(_01787_),
    .A2(_01798_),
    .B(_01804_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09411_ (.I(_01029_),
    .Z(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09412_ (.I(_01805_),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09413_ (.I(_01797_),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09414_ (.I(_01797_),
    .Z(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09415_ (.A1(\filters.lp ),
    .A2(_01808_),
    .B(_01801_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09416_ (.A1(_01806_),
    .A2(_01807_),
    .B(_01809_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09417_ (.I(_01042_),
    .Z(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09418_ (.I(_01810_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09419_ (.I(_01811_),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09420_ (.I(_01762_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09421_ (.A1(\filters.bp ),
    .A2(_01808_),
    .B(_01813_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09422_ (.A1(_01812_),
    .A2(_01807_),
    .B(_01814_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09423_ (.I(net13),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _09424_ (.I(_01815_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09425_ (.I(_01816_),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09426_ (.I(_01817_),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09427_ (.A1(\filters.hp ),
    .A2(_01808_),
    .B(_01813_),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09428_ (.A1(_01818_),
    .A2(_01807_),
    .B(_01819_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09429_ (.I(net14),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09430_ (.I(_01820_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09431_ (.I(_01821_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09432_ (.I(_01822_),
    .Z(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09433_ (.A1(\filters.mode_vol[7] ),
    .A2(_01808_),
    .B(_01813_),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09434_ (.A1(_01823_),
    .A2(_01807_),
    .B(_01824_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09435_ (.I(_01028_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09436_ (.I(_01825_),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09437_ (.I(_01826_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09438_ (.I(_01827_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09439_ (.I(_01014_),
    .Z(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09440_ (.I(_01829_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09441_ (.I(net3),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _09442_ (.A1(_01792_),
    .A2(net4),
    .A3(_01831_),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09443_ (.A1(_01830_),
    .A2(_01832_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09444_ (.I(_01833_),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09445_ (.I(net5),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09446_ (.I(_01835_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09447_ (.A1(net4),
    .A2(net3),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09448_ (.I(_01837_),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09449_ (.A1(_01836_),
    .A2(_01830_),
    .A3(_01838_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09450_ (.I(_01839_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09451_ (.A1(\channels.ctrl_reg2[0] ),
    .A2(_01834_),
    .B1(_01840_),
    .B2(\channels.freq3[8] ),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09452_ (.I(_01835_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09453_ (.I(_01793_),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09454_ (.A1(_01842_),
    .A2(_01843_),
    .A3(_01838_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09455_ (.I(_01844_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09456_ (.I(_01792_),
    .Z(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09457_ (.I(net2),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09458_ (.A1(_01847_),
    .A2(net1),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09459_ (.I(_01848_),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09460_ (.A1(_01012_),
    .A2(_01831_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09461_ (.I(_01850_),
    .Z(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09462_ (.A1(_01846_),
    .A2(_01849_),
    .A3(_01851_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09463_ (.I(_01852_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09464_ (.A1(\channels.atk_dec2[0] ),
    .A2(_01845_),
    .B1(_01853_),
    .B2(\channels.pw3[8] ),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09465_ (.I(_01015_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09466_ (.A1(_01849_),
    .A2(_01832_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09467_ (.I(_01856_),
    .Z(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09468_ (.I(_01013_),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09469_ (.I(_01858_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09470_ (.A1(_01846_),
    .A2(_01859_),
    .A3(_01848_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09471_ (.A1(_01847_),
    .A2(net1),
    .Z(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09472_ (.A1(_01792_),
    .A2(_01858_),
    .A3(_01861_),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09473_ (.A1(\filters.cutoff_lut[6] ),
    .A2(_01860_),
    .B1(_01862_),
    .B2(\filters.cutoff_lut[9] ),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09474_ (.I(net5),
    .Z(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09475_ (.I(_01850_),
    .Z(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09476_ (.A1(_01864_),
    .A2(_01843_),
    .A3(_01865_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09477_ (.A1(_01864_),
    .A2(_01858_),
    .A3(_01843_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09478_ (.A1(\channels.freq1[0] ),
    .A2(_01866_),
    .B1(_01867_),
    .B2(\channels.ctrl_reg1[0] ),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09479_ (.A1(_01858_),
    .A2(_01794_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09480_ (.A1(_01861_),
    .A2(_01832_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09481_ (.I(_01870_),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09482_ (.A1(\channels.sus_rel3[0] ),
    .A2(_01869_),
    .B1(_01871_),
    .B2(\channels.pw2[8] ),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09483_ (.A1(_01863_),
    .A2(_01868_),
    .A3(_01872_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09484_ (.A1(_01758_),
    .A2(_01855_),
    .B1(_01857_),
    .B2(\channels.pw2[0] ),
    .C(_01873_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09485_ (.A1(_01846_),
    .A2(_01829_),
    .A3(_01865_),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09486_ (.I(_01875_),
    .Z(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09487_ (.A1(_01836_),
    .A2(_01848_),
    .A3(_01838_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09488_ (.I(_01877_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09489_ (.I(_01861_),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09490_ (.A1(_01836_),
    .A2(_01879_),
    .A3(_01838_),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09491_ (.I(_01880_),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09492_ (.A1(\channels.atk_dec3[0] ),
    .A2(_01876_),
    .B1(_01878_),
    .B2(\channels.sus_rel2[0] ),
    .C1(_01881_),
    .C2(\channels.freq3[0] ),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09493_ (.A1(_01841_),
    .A2(_01854_),
    .A3(_01874_),
    .A4(_01882_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09494_ (.I(net6),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09495_ (.I(_01884_),
    .Z(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09496_ (.A1(_01794_),
    .A2(_01837_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09497_ (.I(_01886_),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09498_ (.A1(\channels.ch3_env[0] ),
    .A2(_01887_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09499_ (.A1(_01842_),
    .A2(_01859_),
    .A3(_01830_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09500_ (.I(_01889_),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09501_ (.A1(_01846_),
    .A2(_01879_),
    .A3(_01851_),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09502_ (.I(_01891_),
    .Z(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09503_ (.A1(\channels.freq2[0] ),
    .A2(_01890_),
    .B1(_01892_),
    .B2(\channels.ctrl_reg3[0] ),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09504_ (.A1(_01864_),
    .A2(_01879_),
    .A3(_01865_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09505_ (.I(_01894_),
    .Z(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09506_ (.A1(_01864_),
    .A2(_01848_),
    .A3(_01865_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09507_ (.I(_01896_),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09508_ (.A1(\channels.pw1[0] ),
    .A2(_01895_),
    .B1(_01897_),
    .B2(\channels.freq1[8] ),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09509_ (.A1(_01885_),
    .A2(_01888_),
    .A3(_01893_),
    .A4(_01898_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09510_ (.A1(_01842_),
    .A2(_01829_),
    .A3(_01851_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09511_ (.I(_01900_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09512_ (.A1(_01843_),
    .A2(_01832_),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09513_ (.I(_01902_),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09514_ (.A1(\channels.pw1[8] ),
    .A2(_01901_),
    .B1(_01903_),
    .B2(\channels.freq2[8] ),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09515_ (.I(_01795_),
    .Z(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09516_ (.A1(_01794_),
    .A2(_01851_),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09517_ (.I(_01906_),
    .Z(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09518_ (.A1(\filters.mode_vol[0] ),
    .A2(_01905_),
    .B1(_01907_),
    .B2(\channels.pw3[0] ),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09519_ (.A1(_01836_),
    .A2(_01859_),
    .A3(_01879_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09520_ (.I(_01909_),
    .Z(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09521_ (.A1(_01842_),
    .A2(_01859_),
    .A3(_01849_),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09522_ (.I(_01911_),
    .Z(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09523_ (.A1(\channels.sus_rel1[0] ),
    .A2(_01910_),
    .B1(_01912_),
    .B2(\channels.atk_dec1[0] ),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09524_ (.A1(_01835_),
    .A2(net4),
    .A3(_01831_),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09525_ (.A1(_01830_),
    .A2(_01914_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09526_ (.I(_01915_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09527_ (.A1(_01849_),
    .A2(_01914_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09528_ (.A1(\channels.sample3[4] ),
    .A2(_01916_),
    .B1(_01917_),
    .B2(\clk_trg[0] ),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09529_ (.A1(_01904_),
    .A2(_01908_),
    .A3(_01913_),
    .A4(_01918_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09530_ (.I(_01884_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09531_ (.I(_01920_),
    .Z(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09532_ (.A1(_01883_),
    .A2(_01899_),
    .A3(_01919_),
    .B1(net21),
    .B2(_01921_),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09533_ (.A1(_01828_),
    .A2(_01922_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09534_ (.A1(\channels.ctrl_reg2[1] ),
    .A2(_01834_),
    .B1(_01840_),
    .B2(\channels.freq3[9] ),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09535_ (.A1(\channels.atk_dec2[1] ),
    .A2(_01845_),
    .B1(_01853_),
    .B2(\channels.pw3[9] ),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09536_ (.A1(\filters.cutoff_lut[7] ),
    .A2(_01860_),
    .B1(_01862_),
    .B2(\filters.cutoff_lut[10] ),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09537_ (.A1(\channels.freq1[1] ),
    .A2(_01866_),
    .B1(_01867_),
    .B2(\channels.ctrl_reg1[1] ),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09538_ (.A1(\channels.sus_rel3[1] ),
    .A2(_01869_),
    .B1(_01870_),
    .B2(\channels.pw2[9] ),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09539_ (.A1(_01925_),
    .A2(_01926_),
    .A3(_01927_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09540_ (.A1(_01772_),
    .A2(_01855_),
    .B1(_01857_),
    .B2(\channels.pw2[1] ),
    .C(_01928_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09541_ (.A1(\channels.atk_dec3[1] ),
    .A2(_01876_),
    .B1(_01878_),
    .B2(\channels.sus_rel2[1] ),
    .C1(_01881_),
    .C2(\channels.freq3[1] ),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09542_ (.A1(_01923_),
    .A2(_01924_),
    .A3(_01929_),
    .A4(_01930_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09543_ (.A1(\channels.ch3_env[1] ),
    .A2(_01887_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09544_ (.A1(\channels.freq2[1] ),
    .A2(_01890_),
    .B1(_01892_),
    .B2(\channels.ctrl_reg3[1] ),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09545_ (.A1(\channels.pw1[1] ),
    .A2(_01895_),
    .B1(_01897_),
    .B2(\channels.freq1[9] ),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09546_ (.A1(_01885_),
    .A2(_01932_),
    .A3(_01933_),
    .A4(_01934_),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09547_ (.A1(\channels.pw1[9] ),
    .A2(_01901_),
    .B1(_01903_),
    .B2(\channels.freq2[9] ),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09548_ (.A1(\filters.mode_vol[1] ),
    .A2(_01796_),
    .B1(_01907_),
    .B2(\channels.pw3[1] ),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09549_ (.A1(\channels.sus_rel1[1] ),
    .A2(_01910_),
    .B1(_01912_),
    .B2(\channels.atk_dec1[1] ),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09550_ (.I(\channels.sample3[5] ),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09551_ (.A1(_01939_),
    .A2(_01916_),
    .B1(_01917_),
    .B2(\clk_trg[1] ),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09552_ (.A1(_01936_),
    .A2(_01937_),
    .A3(_01938_),
    .A4(_01940_),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09553_ (.A1(_01931_),
    .A2(_01935_),
    .A3(_01941_),
    .B1(net22),
    .B2(_01921_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09554_ (.A1(_01828_),
    .A2(_01942_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09555_ (.I(_01052_),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09556_ (.I(_01943_),
    .Z(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09557_ (.I(_01944_),
    .Z(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09558_ (.I(_01884_),
    .Z(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09559_ (.A1(\channels.ctrl_reg3[2] ),
    .A2(_01892_),
    .B1(_01871_),
    .B2(\channels.pw2[10] ),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09560_ (.I(_01877_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09561_ (.I(_01880_),
    .Z(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09562_ (.A1(\channels.sus_rel2[2] ),
    .A2(_01948_),
    .B1(_01949_),
    .B2(\channels.freq3[2] ),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09563_ (.I(_01916_),
    .Z(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09564_ (.A1(_01783_),
    .A2(_01015_),
    .B1(_01795_),
    .B2(\filters.mode_vol[2] ),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09565_ (.I(_01867_),
    .Z(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09566_ (.A1(\channels.pw1[10] ),
    .A2(_01900_),
    .B1(_01953_),
    .B2(\channels.ctrl_reg1[2] ),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09567_ (.I(_01869_),
    .Z(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09568_ (.A1(\filters.cutoff_lut[8] ),
    .A2(_01860_),
    .B1(_01955_),
    .B2(\channels.sus_rel3[2] ),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09569_ (.A1(_01952_),
    .A2(_01954_),
    .A3(_01956_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09570_ (.A1(\channels.sus_rel1[2] ),
    .A2(_01910_),
    .B1(_01951_),
    .B2(\channels.sample3[6] ),
    .C(_01957_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09571_ (.A1(_01947_),
    .A2(_01950_),
    .A3(_01958_),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09572_ (.I(_01911_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09573_ (.A1(\channels.atk_dec1[2] ),
    .A2(_01960_),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09574_ (.A1(\channels.pw1[2] ),
    .A2(_01894_),
    .B1(_01902_),
    .B2(\channels.freq2[10] ),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09575_ (.A1(\channels.ctrl_reg2[2] ),
    .A2(_01833_),
    .B1(_01889_),
    .B2(\channels.freq2[2] ),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09576_ (.A1(_01962_),
    .A2(_01963_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09577_ (.A1(\channels.pw3[10] ),
    .A2(_01853_),
    .B1(_01857_),
    .B2(\channels.pw2[2] ),
    .C(_01964_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09578_ (.I(_01866_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09579_ (.A1(\channels.ch3_env[2] ),
    .A2(_01886_),
    .B1(_01896_),
    .B2(\channels.freq1[10] ),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09580_ (.I(_01862_),
    .Z(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09581_ (.A1(\filters.cutoff_lut[11] ),
    .A2(_01968_),
    .B1(_01875_),
    .B2(\channels.atk_dec3[2] ),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09582_ (.A1(\channels.atk_dec2[2] ),
    .A2(_01844_),
    .B1(_01906_),
    .B2(\channels.pw3[2] ),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09583_ (.A1(_01967_),
    .A2(_01969_),
    .A3(_01970_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09584_ (.A1(\channels.freq1[2] ),
    .A2(_01966_),
    .B1(_01840_),
    .B2(\channels.freq3[10] ),
    .C(_01971_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09585_ (.A1(_01885_),
    .A2(_01961_),
    .A3(_01965_),
    .A4(_01972_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09586_ (.A1(_01946_),
    .A2(net23),
    .B1(_01959_),
    .B2(_01973_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09587_ (.A1(_01945_),
    .A2(_01974_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09588_ (.I(_01955_),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09589_ (.I(_01909_),
    .Z(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09590_ (.A1(\channels.sus_rel3[3] ),
    .A2(_01975_),
    .B1(_01976_),
    .B2(\channels.sus_rel1[3] ),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09591_ (.I(_01844_),
    .Z(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09592_ (.A1(\filters.res_filt[3] ),
    .A2(_01855_),
    .B1(_01903_),
    .B2(\channels.freq2[11] ),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09593_ (.A1(\filters.mode_vol[3] ),
    .A2(_01796_),
    .B1(_01877_),
    .B2(\channels.sus_rel2[3] ),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09594_ (.A1(\channels.ch3_env[3] ),
    .A2(_01887_),
    .B1(_01895_),
    .B2(\channels.pw1[3] ),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09595_ (.I(_01896_),
    .Z(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09596_ (.A1(\channels.pw3[11] ),
    .A2(_01852_),
    .B1(_01982_),
    .B2(\channels.freq1[11] ),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09597_ (.A1(_01979_),
    .A2(_01980_),
    .A3(_01981_),
    .A4(_01983_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09598_ (.A1(\channels.atk_dec2[3] ),
    .A2(_01978_),
    .B(_01984_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09599_ (.I(_01833_),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09600_ (.A1(\channels.pw1[11] ),
    .A2(_01901_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09601_ (.A1(\channels.freq3[3] ),
    .A2(_01880_),
    .B1(_01889_),
    .B2(\channels.freq2[3] ),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09602_ (.I(\channels.sample3[7] ),
    .Z(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09603_ (.A1(\channels.ctrl_reg1[3] ),
    .A2(_01953_),
    .B1(_01915_),
    .B2(_01989_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09604_ (.A1(_01884_),
    .A2(_01987_),
    .A3(_01988_),
    .A4(_01990_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09605_ (.A1(\channels.ctrl_reg2[3] ),
    .A2(_01986_),
    .B1(_01892_),
    .B2(\channels.ctrl_reg3[3] ),
    .C(_01991_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09606_ (.A1(\channels.pw2[3] ),
    .A2(_01856_),
    .B1(_01911_),
    .B2(\channels.atk_dec1[3] ),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09607_ (.A1(\channels.atk_dec3[3] ),
    .A2(_01876_),
    .B1(_01906_),
    .B2(\channels.pw3[3] ),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09608_ (.A1(\filters.cutoff_lut[12] ),
    .A2(_01968_),
    .B1(_01866_),
    .B2(\channels.freq1[3] ),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09609_ (.A1(_01993_),
    .A2(_01994_),
    .A3(_01995_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09610_ (.A1(\channels.freq3[11] ),
    .A2(_01840_),
    .B1(_01871_),
    .B2(\channels.pw2[11] ),
    .C(_01996_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09611_ (.A1(_01977_),
    .A2(_01985_),
    .A3(_01992_),
    .A4(_01997_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09612_ (.A1(_01921_),
    .A2(net24),
    .B(_01998_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09613_ (.A1(_01945_),
    .A2(_01999_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09614_ (.I(_01968_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09615_ (.A1(\filters.cutoff_lut[13] ),
    .A2(_02000_),
    .ZN(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09616_ (.A1(\channels.sus_rel3[4] ),
    .A2(_01975_),
    .B1(_01897_),
    .B2(\channels.freq1[12] ),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09617_ (.I(_01875_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09618_ (.I(_01839_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09619_ (.A1(\channels.atk_dec3[4] ),
    .A2(_02003_),
    .B1(_02004_),
    .B2(\channels.freq3[12] ),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09620_ (.A1(_01885_),
    .A2(_02001_),
    .A3(_02002_),
    .A4(_02005_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09621_ (.A1(\channels.ctrl_reg2[4] ),
    .A2(_01986_),
    .B1(_01978_),
    .B2(\channels.atk_dec2[4] ),
    .C(_02006_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09622_ (.I(_01856_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09623_ (.I(_01902_),
    .Z(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09624_ (.A1(\channels.pw2[4] ),
    .A2(_02008_),
    .B1(_02009_),
    .B2(\channels.freq2[12] ),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09625_ (.I(_01891_),
    .Z(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09626_ (.A1(\channels.freq3[4] ),
    .A2(_01949_),
    .B1(_02011_),
    .B2(\channels.ctrl_reg3[4] ),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09627_ (.I(_01889_),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09628_ (.A1(\channels.sus_rel2[4] ),
    .A2(_01948_),
    .B1(_02013_),
    .B2(\channels.freq2[4] ),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09629_ (.I(_01894_),
    .Z(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09630_ (.I(_01953_),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09631_ (.A1(\channels.pw1[4] ),
    .A2(_02015_),
    .B1(_02016_),
    .B2(\channels.ctrl_reg1[4] ),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09632_ (.A1(_02010_),
    .A2(_02012_),
    .A3(_02014_),
    .A4(_02017_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09633_ (.I(_01855_),
    .Z(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09634_ (.A1(\filters.res_filt[4] ),
    .A2(_02019_),
    .B1(_01951_),
    .B2(\channels.sample3[8] ),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09635_ (.I(_01887_),
    .Z(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09636_ (.A1(\channels.ch3_env[4] ),
    .A2(_02021_),
    .B1(_01960_),
    .B2(\channels.atk_dec1[4] ),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09637_ (.I(_01966_),
    .Z(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09638_ (.I(_01906_),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09639_ (.A1(\channels.freq1[4] ),
    .A2(_02023_),
    .B1(_02024_),
    .B2(\channels.pw3[4] ),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09640_ (.A1(\filters.lp ),
    .A2(_01905_),
    .B1(_01976_),
    .B2(\channels.sus_rel1[4] ),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09641_ (.A1(_02020_),
    .A2(_02022_),
    .A3(_02025_),
    .A4(_02026_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09642_ (.A1(_02018_),
    .A2(_02027_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09643_ (.A1(_01946_),
    .A2(net25),
    .B(_01813_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09644_ (.A1(_02007_),
    .A2(_02028_),
    .B(_02029_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09645_ (.A1(\filters.cutoff_lut[14] ),
    .A2(_02000_),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09646_ (.A1(\channels.sus_rel3[5] ),
    .A2(_01975_),
    .B1(_01982_),
    .B2(\channels.freq1[13] ),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09647_ (.A1(\channels.atk_dec3[5] ),
    .A2(_02003_),
    .B1(_02004_),
    .B2(\channels.freq3[13] ),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09648_ (.A1(_01920_),
    .A2(_02030_),
    .A3(_02031_),
    .A4(_02032_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09649_ (.A1(\channels.ctrl_reg2[5] ),
    .A2(_01986_),
    .B1(_01978_),
    .B2(\channels.atk_dec2[5] ),
    .C(_02033_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09650_ (.A1(\channels.pw2[5] ),
    .A2(_02008_),
    .B1(_02009_),
    .B2(\channels.freq2[13] ),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09651_ (.A1(\channels.freq3[5] ),
    .A2(_01881_),
    .B1(_02011_),
    .B2(\channels.ctrl_reg3[5] ),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09652_ (.A1(\channels.sus_rel2[5] ),
    .A2(_01948_),
    .B1(_02013_),
    .B2(\channels.freq2[5] ),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09653_ (.A1(\channels.pw1[5] ),
    .A2(_02015_),
    .B1(_02016_),
    .B2(\channels.ctrl_reg1[5] ),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09654_ (.A1(_02035_),
    .A2(_02036_),
    .A3(_02037_),
    .A4(_02038_),
    .ZN(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09655_ (.I(\channels.sample3[9] ),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09656_ (.A1(\filters.res_filt[5] ),
    .A2(_02019_),
    .B1(_01951_),
    .B2(_02040_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09657_ (.A1(\channels.ch3_env[5] ),
    .A2(_02021_),
    .B1(_01960_),
    .B2(\channels.atk_dec1[5] ),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09658_ (.A1(\channels.freq1[5] ),
    .A2(_02023_),
    .B1(_02024_),
    .B2(\channels.pw3[5] ),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09659_ (.A1(\filters.bp ),
    .A2(_01905_),
    .B1(_01976_),
    .B2(\channels.sus_rel1[5] ),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09660_ (.A1(_02041_),
    .A2(_02042_),
    .A3(_02043_),
    .A4(_02044_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09661_ (.A1(_02039_),
    .A2(_02045_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09662_ (.I(_01761_),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09663_ (.I(_02047_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09664_ (.A1(_01946_),
    .A2(net26),
    .B(_02048_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09665_ (.A1(_02034_),
    .A2(_02046_),
    .B(_02049_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09666_ (.A1(\filters.cutoff_lut[15] ),
    .A2(_02000_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09667_ (.A1(\channels.sus_rel3[6] ),
    .A2(_01955_),
    .B1(_01982_),
    .B2(\channels.freq1[14] ),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09668_ (.A1(\channels.atk_dec3[6] ),
    .A2(_02003_),
    .B1(_02004_),
    .B2(\channels.freq3[14] ),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09669_ (.A1(_01920_),
    .A2(_02050_),
    .A3(_02051_),
    .A4(_02052_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09670_ (.A1(\channels.ctrl_reg2[6] ),
    .A2(_01986_),
    .B1(_01978_),
    .B2(\channels.atk_dec2[6] ),
    .C(_02053_),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09671_ (.A1(\channels.pw2[6] ),
    .A2(_01857_),
    .B1(_02009_),
    .B2(\channels.freq2[14] ),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09672_ (.A1(\channels.freq3[6] ),
    .A2(_01881_),
    .B1(_02011_),
    .B2(\channels.ctrl_reg3[6] ),
    .ZN(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09673_ (.A1(\channels.sus_rel2[6] ),
    .A2(_01878_),
    .B1(_01890_),
    .B2(\channels.freq2[6] ),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09674_ (.A1(\channels.pw1[6] ),
    .A2(_01895_),
    .B1(_02016_),
    .B2(\channels.ctrl_reg1[6] ),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09675_ (.A1(_02055_),
    .A2(_02056_),
    .A3(_02057_),
    .A4(_02058_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09676_ (.A1(\filters.res_filt[6] ),
    .A2(_02019_),
    .B1(_01951_),
    .B2(\channels.sample3[10] ),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09677_ (.A1(\channels.ch3_env[6] ),
    .A2(_02021_),
    .B1(_01960_),
    .B2(\channels.atk_dec1[6] ),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09678_ (.A1(\channels.freq1[6] ),
    .A2(_02023_),
    .B1(_02024_),
    .B2(\channels.pw3[6] ),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09679_ (.A1(\filters.hp ),
    .A2(_01905_),
    .B1(_01910_),
    .B2(\channels.sus_rel1[6] ),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09680_ (.A1(_02060_),
    .A2(_02061_),
    .A3(_02062_),
    .A4(_02063_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09681_ (.A1(_02059_),
    .A2(_02064_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09682_ (.A1(_01946_),
    .A2(net27),
    .B(_02048_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09683_ (.A1(_02054_),
    .A2(_02065_),
    .B(_02066_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09684_ (.A1(\filters.mode_vol[7] ),
    .A2(_01796_),
    .B1(_02004_),
    .B2(\channels.freq3[15] ),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09685_ (.I(\channels.sample3[11] ),
    .Z(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09686_ (.A1(\channels.ctrl_reg2[7] ),
    .A2(_01834_),
    .B1(_01916_),
    .B2(_02068_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09687_ (.A1(\channels.atk_dec1[7] ),
    .A2(_01912_),
    .B(_01917_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09688_ (.A1(_01920_),
    .A2(_02067_),
    .A3(_02069_),
    .A4(_02070_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09689_ (.A1(\channels.ch3_env[7] ),
    .A2(_02021_),
    .B1(_01976_),
    .B2(\channels.sus_rel1[7] ),
    .C(_02071_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09690_ (.A1(\channels.freq1[7] ),
    .A2(_01966_),
    .B1(_01948_),
    .B2(\channels.sus_rel2[7] ),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09691_ (.A1(\channels.atk_dec3[7] ),
    .A2(_02003_),
    .B1(_02013_),
    .B2(\channels.freq2[7] ),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09692_ (.A1(\channels.freq2[15] ),
    .A2(_02009_),
    .B1(_01897_),
    .B2(\channels.freq1[15] ),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09693_ (.A1(\channels.atk_dec2[7] ),
    .A2(_01845_),
    .B1(_01949_),
    .B2(\channels.freq3[7] ),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09694_ (.A1(_02073_),
    .A2(_02074_),
    .A3(_02075_),
    .A4(_02076_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09695_ (.A1(\channels.ctrl_reg3[7] ),
    .A2(_02011_),
    .B1(_02016_),
    .B2(\channels.ctrl_reg1[7] ),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09696_ (.A1(\filters.cutoff_lut[16] ),
    .A2(_02000_),
    .B1(_01975_),
    .B2(\channels.sus_rel3[7] ),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09697_ (.A1(\filters.res_filt[7] ),
    .A2(_02019_),
    .B1(_01907_),
    .B2(\channels.pw3[7] ),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09698_ (.A1(\channels.pw1[7] ),
    .A2(_02015_),
    .B1(_02008_),
    .B2(\channels.pw2[7] ),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09699_ (.A1(_02078_),
    .A2(_02079_),
    .A3(_02080_),
    .A4(_02081_),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09700_ (.A1(_02077_),
    .A2(_02082_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09701_ (.A1(net28),
    .A2(_01921_),
    .B(_02048_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09702_ (.A1(_02072_),
    .A2(_02083_),
    .B(_02084_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09703_ (.A1(_01791_),
    .A2(_01982_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09704_ (.I(_02085_),
    .Z(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09705_ (.I(_02085_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09706_ (.A1(\channels.freq1[8] ),
    .A2(_02087_),
    .B(_02048_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09707_ (.A1(_01752_),
    .A2(_02086_),
    .B(_02088_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09708_ (.I(_02047_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09709_ (.A1(\channels.freq1[9] ),
    .A2(_02087_),
    .B(_02089_),
    .ZN(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09710_ (.A1(_01767_),
    .A2(_02086_),
    .B(_02090_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09711_ (.A1(\channels.freq1[10] ),
    .A2(_02087_),
    .B(_02089_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09712_ (.A1(_01777_),
    .A2(_02086_),
    .B(_02091_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09713_ (.A1(\channels.freq1[11] ),
    .A2(_02087_),
    .B(_02089_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09714_ (.A1(_01787_),
    .A2(_02086_),
    .B(_02092_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09715_ (.I(_02085_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09716_ (.I(_02085_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09717_ (.A1(\channels.freq1[12] ),
    .A2(_02094_),
    .B(_02089_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09718_ (.A1(_01806_),
    .A2(_02093_),
    .B(_02095_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09719_ (.I(_02047_),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09720_ (.A1(\channels.freq1[13] ),
    .A2(_02094_),
    .B(_02096_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09721_ (.A1(_01812_),
    .A2(_02093_),
    .B(_02097_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09722_ (.A1(\channels.freq1[14] ),
    .A2(_02094_),
    .B(_02096_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09723_ (.A1(_01818_),
    .A2(_02093_),
    .B(_02098_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09724_ (.A1(\channels.freq1[15] ),
    .A2(_02094_),
    .B(_02096_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09725_ (.A1(_01823_),
    .A2(_02093_),
    .B(_02099_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09726_ (.I(_01790_),
    .Z(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09727_ (.A1(_02100_),
    .A2(_01901_),
    .Z(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09728_ (.I(_02101_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09729_ (.I(_02101_),
    .Z(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09730_ (.A1(\channels.pw1[8] ),
    .A2(_02103_),
    .B(_02096_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09731_ (.A1(_01752_),
    .A2(_02102_),
    .B(_02104_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09732_ (.I(_02047_),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09733_ (.A1(\channels.pw1[9] ),
    .A2(_02103_),
    .B(_02105_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09734_ (.A1(_01767_),
    .A2(_02102_),
    .B(_02106_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09735_ (.A1(\channels.pw1[10] ),
    .A2(_02103_),
    .B(_02105_),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09736_ (.A1(_01777_),
    .A2(_02102_),
    .B(_02107_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09737_ (.A1(\channels.pw1[11] ),
    .A2(_02103_),
    .B(_02105_),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09738_ (.A1(_01787_),
    .A2(_02102_),
    .B(_02108_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09739_ (.I(_01749_),
    .Z(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09740_ (.I(_02109_),
    .Z(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09741_ (.A1(_01791_),
    .A2(_01953_),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09742_ (.I(_02111_),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09743_ (.I(_02111_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09744_ (.A1(\channels.ctrl_reg1[0] ),
    .A2(_02113_),
    .B(_02105_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09745_ (.A1(_02110_),
    .A2(_02112_),
    .B(_02114_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09746_ (.I(_01766_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09747_ (.I(_01760_),
    .Z(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09748_ (.I(_02116_),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09749_ (.I(_02117_),
    .Z(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09750_ (.A1(\channels.ctrl_reg1[1] ),
    .A2(_02113_),
    .B(_02118_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09751_ (.A1(_02115_),
    .A2(_02112_),
    .B(_02119_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09752_ (.I(_01776_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09753_ (.A1(\channels.ctrl_reg1[2] ),
    .A2(_02113_),
    .B(_02118_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09754_ (.A1(_02120_),
    .A2(_02112_),
    .B(_02121_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09755_ (.I(_01786_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09756_ (.A1(\channels.ctrl_reg1[3] ),
    .A2(_02113_),
    .B(_02118_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09757_ (.A1(_02122_),
    .A2(_02112_),
    .B(_02123_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09758_ (.I(_02111_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09759_ (.I(_02111_),
    .Z(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09760_ (.A1(\channels.ctrl_reg1[4] ),
    .A2(_02125_),
    .B(_02118_),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09761_ (.A1(_01806_),
    .A2(_02124_),
    .B(_02126_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09762_ (.I(_02117_),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09763_ (.A1(\channels.ctrl_reg1[5] ),
    .A2(_02125_),
    .B(_02127_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09764_ (.A1(_01812_),
    .A2(_02124_),
    .B(_02128_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09765_ (.A1(\channels.ctrl_reg1[6] ),
    .A2(_02125_),
    .B(_02127_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09766_ (.A1(_01818_),
    .A2(_02124_),
    .B(_02129_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09767_ (.A1(\channels.ctrl_reg1[7] ),
    .A2(_02125_),
    .B(_02127_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09768_ (.A1(_01823_),
    .A2(_02124_),
    .B(_02130_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09769_ (.A1(_01791_),
    .A2(_01912_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09770_ (.I(_02131_),
    .Z(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09771_ (.I(_02131_),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09772_ (.A1(\channels.atk_dec1[0] ),
    .A2(_02133_),
    .B(_02127_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09773_ (.A1(_02110_),
    .A2(_02132_),
    .B(_02134_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09774_ (.I(_02117_),
    .Z(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09775_ (.A1(\channels.atk_dec1[1] ),
    .A2(_02133_),
    .B(_02135_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09776_ (.A1(_02115_),
    .A2(_02132_),
    .B(_02136_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09777_ (.A1(\channels.atk_dec1[2] ),
    .A2(_02133_),
    .B(_02135_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09778_ (.A1(_02120_),
    .A2(_02132_),
    .B(_02137_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09779_ (.A1(\channels.atk_dec1[3] ),
    .A2(_02133_),
    .B(_02135_),
    .ZN(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09780_ (.A1(_02122_),
    .A2(_02132_),
    .B(_02138_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09781_ (.I(_02131_),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09782_ (.I(_02131_),
    .Z(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09783_ (.A1(\channels.atk_dec1[4] ),
    .A2(_02140_),
    .B(_02135_),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09784_ (.A1(_01806_),
    .A2(_02139_),
    .B(_02141_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09785_ (.I(_02117_),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09786_ (.A1(\channels.atk_dec1[5] ),
    .A2(_02140_),
    .B(_02142_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09787_ (.A1(_01812_),
    .A2(_02139_),
    .B(_02143_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09788_ (.A1(\channels.atk_dec1[6] ),
    .A2(_02140_),
    .B(_02142_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09789_ (.A1(_01818_),
    .A2(_02139_),
    .B(_02144_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09790_ (.A1(\channels.atk_dec1[7] ),
    .A2(_02140_),
    .B(_02142_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09791_ (.A1(_01823_),
    .A2(_02139_),
    .B(_02145_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09792_ (.I(_01790_),
    .Z(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09793_ (.A1(_02146_),
    .A2(_01909_),
    .Z(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09794_ (.I(_02147_),
    .Z(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09795_ (.I(_02147_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09796_ (.A1(\channels.sus_rel1[0] ),
    .A2(_02149_),
    .B(_02142_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09797_ (.A1(_02110_),
    .A2(_02148_),
    .B(_02150_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09798_ (.I(_02116_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09799_ (.I(_02151_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09800_ (.A1(\channels.sus_rel1[1] ),
    .A2(_02149_),
    .B(_02152_),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09801_ (.A1(_02115_),
    .A2(_02148_),
    .B(_02153_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09802_ (.A1(\channels.sus_rel1[2] ),
    .A2(_02149_),
    .B(_02152_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09803_ (.A1(_02120_),
    .A2(_02148_),
    .B(_02154_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09804_ (.A1(\channels.sus_rel1[3] ),
    .A2(_02149_),
    .B(_02152_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09805_ (.A1(_02122_),
    .A2(_02148_),
    .B(_02155_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09806_ (.I(_01805_),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09807_ (.I(_02147_),
    .Z(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09808_ (.I(_02147_),
    .Z(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09809_ (.A1(\channels.sus_rel1[4] ),
    .A2(_02158_),
    .B(_02152_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09810_ (.A1(_02156_),
    .A2(_02157_),
    .B(_02159_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09811_ (.I(_01810_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09812_ (.I(_02160_),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09813_ (.I(_02151_),
    .Z(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09814_ (.A1(\channels.sus_rel1[5] ),
    .A2(_02158_),
    .B(_02162_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09815_ (.A1(_02161_),
    .A2(_02157_),
    .B(_02163_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09816_ (.I(_01817_),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09817_ (.A1(\channels.sus_rel1[6] ),
    .A2(_02158_),
    .B(_02162_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09818_ (.A1(_02164_),
    .A2(_02157_),
    .B(_02165_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09819_ (.I(_01822_),
    .Z(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09820_ (.A1(\channels.sus_rel1[7] ),
    .A2(_02158_),
    .B(_02162_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09821_ (.A1(_02166_),
    .A2(_02157_),
    .B(_02167_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09822_ (.A1(_02146_),
    .A2(_01903_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09823_ (.I(_02168_),
    .Z(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09824_ (.I(_02168_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09825_ (.A1(\channels.freq2[8] ),
    .A2(_02170_),
    .B(_02162_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09826_ (.A1(_02110_),
    .A2(_02169_),
    .B(_02171_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09827_ (.I(_02151_),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09828_ (.A1(\channels.freq2[9] ),
    .A2(_02170_),
    .B(_02172_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09829_ (.A1(_02115_),
    .A2(_02169_),
    .B(_02173_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09830_ (.A1(\channels.freq2[10] ),
    .A2(_02170_),
    .B(_02172_),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09831_ (.A1(_02120_),
    .A2(_02169_),
    .B(_02174_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09832_ (.A1(\channels.freq2[11] ),
    .A2(_02170_),
    .B(_02172_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09833_ (.A1(_02122_),
    .A2(_02169_),
    .B(_02175_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09834_ (.I(_02168_),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09835_ (.I(_02168_),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09836_ (.A1(\channels.freq2[12] ),
    .A2(_02177_),
    .B(_02172_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09837_ (.A1(_02156_),
    .A2(_02176_),
    .B(_02178_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09838_ (.I(_02151_),
    .Z(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09839_ (.A1(\channels.freq2[13] ),
    .A2(_02177_),
    .B(_02179_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09840_ (.A1(_02161_),
    .A2(_02176_),
    .B(_02180_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09841_ (.A1(\channels.freq2[14] ),
    .A2(_02177_),
    .B(_02179_),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09842_ (.A1(_02164_),
    .A2(_02176_),
    .B(_02181_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09843_ (.A1(\channels.freq2[15] ),
    .A2(_02177_),
    .B(_02179_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09844_ (.A1(_02166_),
    .A2(_02176_),
    .B(_02182_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09845_ (.I(_02109_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09846_ (.A1(_02100_),
    .A2(_01871_),
    .Z(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09847_ (.I(_02184_),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09848_ (.I(_02184_),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09849_ (.A1(\channels.pw2[8] ),
    .A2(_02186_),
    .B(_02179_),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09850_ (.A1(_02183_),
    .A2(_02185_),
    .B(_02187_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09851_ (.I(_01765_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09852_ (.I(_02188_),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09853_ (.I(_02116_),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09854_ (.I(_02190_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09855_ (.A1(\channels.pw2[9] ),
    .A2(_02186_),
    .B(_02191_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09856_ (.A1(_02189_),
    .A2(_02185_),
    .B(_02192_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09857_ (.I(_01775_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09858_ (.I(_02193_),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09859_ (.A1(\channels.pw2[10] ),
    .A2(_02186_),
    .B(_02191_),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09860_ (.A1(_02194_),
    .A2(_02185_),
    .B(_02195_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09861_ (.I(_01786_),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09862_ (.A1(\channels.pw2[11] ),
    .A2(_02186_),
    .B(_02191_),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09863_ (.A1(_02196_),
    .A2(_02185_),
    .B(_02197_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09864_ (.A1(_02146_),
    .A2(_01834_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09865_ (.I(_02198_),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09866_ (.I(_02198_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09867_ (.A1(\channels.ctrl_reg2[0] ),
    .A2(_02200_),
    .B(_02191_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09868_ (.A1(_02183_),
    .A2(_02199_),
    .B(_02201_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09869_ (.I(_02190_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09870_ (.A1(\channels.ctrl_reg2[1] ),
    .A2(_02200_),
    .B(_02202_),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09871_ (.A1(_02189_),
    .A2(_02199_),
    .B(_02203_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09872_ (.A1(\channels.ctrl_reg2[2] ),
    .A2(_02200_),
    .B(_02202_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09873_ (.A1(_02194_),
    .A2(_02199_),
    .B(_02204_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09874_ (.A1(\channels.ctrl_reg2[3] ),
    .A2(_02200_),
    .B(_02202_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09875_ (.A1(_02196_),
    .A2(_02199_),
    .B(_02205_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09876_ (.I(_02198_),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09877_ (.I(_02198_),
    .Z(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09878_ (.A1(\channels.ctrl_reg2[4] ),
    .A2(_02207_),
    .B(_02202_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09879_ (.A1(_02156_),
    .A2(_02206_),
    .B(_02208_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09880_ (.I(_02190_),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09881_ (.A1(\channels.ctrl_reg2[5] ),
    .A2(_02207_),
    .B(_02209_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09882_ (.A1(_02161_),
    .A2(_02206_),
    .B(_02210_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09883_ (.A1(\channels.ctrl_reg2[6] ),
    .A2(_02207_),
    .B(_02209_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09884_ (.A1(_02164_),
    .A2(_02206_),
    .B(_02211_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09885_ (.A1(\channels.ctrl_reg2[7] ),
    .A2(_02207_),
    .B(_02209_),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09886_ (.A1(_02166_),
    .A2(_02206_),
    .B(_02212_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09887_ (.A1(_02146_),
    .A2(_01845_),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09888_ (.I(_02213_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09889_ (.I(_02213_),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09890_ (.A1(\channels.atk_dec2[0] ),
    .A2(_02215_),
    .B(_02209_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09891_ (.A1(_02183_),
    .A2(_02214_),
    .B(_02216_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09892_ (.I(_02190_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09893_ (.A1(\channels.atk_dec2[1] ),
    .A2(_02215_),
    .B(_02217_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09894_ (.A1(_02189_),
    .A2(_02214_),
    .B(_02218_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09895_ (.A1(\channels.atk_dec2[2] ),
    .A2(_02215_),
    .B(_02217_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09896_ (.A1(_02194_),
    .A2(_02214_),
    .B(_02219_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09897_ (.A1(\channels.atk_dec2[3] ),
    .A2(_02215_),
    .B(_02217_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09898_ (.A1(_02196_),
    .A2(_02214_),
    .B(_02220_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09899_ (.I(_02213_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09900_ (.I(_02213_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09901_ (.A1(\channels.atk_dec2[4] ),
    .A2(_02222_),
    .B(_02217_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09902_ (.A1(_02156_),
    .A2(_02221_),
    .B(_02223_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09903_ (.I(_02116_),
    .Z(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09904_ (.I(_02224_),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09905_ (.A1(\channels.atk_dec2[5] ),
    .A2(_02222_),
    .B(_02225_),
    .ZN(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09906_ (.A1(_02161_),
    .A2(_02221_),
    .B(_02226_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09907_ (.A1(\channels.atk_dec2[6] ),
    .A2(_02222_),
    .B(_02225_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09908_ (.A1(_02164_),
    .A2(_02221_),
    .B(_02227_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09909_ (.A1(\channels.atk_dec2[7] ),
    .A2(_02222_),
    .B(_02225_),
    .ZN(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09910_ (.A1(_02166_),
    .A2(_02221_),
    .B(_02228_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09911_ (.I(_01789_),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09912_ (.A1(_02229_),
    .A2(_01878_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09913_ (.I(_02230_),
    .Z(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09914_ (.I(_02230_),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09915_ (.A1(\channels.sus_rel2[0] ),
    .A2(_02232_),
    .B(_02225_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09916_ (.A1(_02183_),
    .A2(_02231_),
    .B(_02233_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09917_ (.I(_02224_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09918_ (.A1(\channels.sus_rel2[1] ),
    .A2(_02232_),
    .B(_02234_),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09919_ (.A1(_02189_),
    .A2(_02231_),
    .B(_02235_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09920_ (.A1(\channels.sus_rel2[2] ),
    .A2(_02232_),
    .B(_02234_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09921_ (.A1(_02194_),
    .A2(_02231_),
    .B(_02236_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09922_ (.A1(\channels.sus_rel2[3] ),
    .A2(_02232_),
    .B(_02234_),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09923_ (.A1(_02196_),
    .A2(_02231_),
    .B(_02237_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09924_ (.I(_01029_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09925_ (.I(_02230_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09926_ (.I(_02230_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09927_ (.A1(\channels.sus_rel2[4] ),
    .A2(_02240_),
    .B(_02234_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09928_ (.A1(_02238_),
    .A2(_02239_),
    .B(_02241_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09929_ (.I(_02160_),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09930_ (.I(_02224_),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09931_ (.A1(\channels.sus_rel2[5] ),
    .A2(_02240_),
    .B(_02243_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09932_ (.A1(_02242_),
    .A2(_02239_),
    .B(_02244_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09933_ (.I(_01817_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09934_ (.A1(\channels.sus_rel2[6] ),
    .A2(_02240_),
    .B(_02243_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09935_ (.A1(_02245_),
    .A2(_02239_),
    .B(_02246_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09936_ (.I(_01822_),
    .Z(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09937_ (.A1(\channels.sus_rel2[7] ),
    .A2(_02240_),
    .B(_02243_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09938_ (.A1(_02247_),
    .A2(_02239_),
    .B(_02248_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09939_ (.I(_02109_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09940_ (.A1(_02229_),
    .A2(_01839_),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09941_ (.I(_02250_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09942_ (.I(_02250_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09943_ (.A1(\channels.freq3[8] ),
    .A2(_02252_),
    .B(_02243_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09944_ (.A1(_02249_),
    .A2(_02251_),
    .B(_02253_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09945_ (.I(_02188_),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09946_ (.I(_02224_),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09947_ (.A1(\channels.freq3[9] ),
    .A2(_02252_),
    .B(_02255_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09948_ (.A1(_02254_),
    .A2(_02251_),
    .B(_02256_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09949_ (.I(_02193_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09950_ (.A1(\channels.freq3[10] ),
    .A2(_02252_),
    .B(_02255_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09951_ (.A1(_02257_),
    .A2(_02251_),
    .B(_02258_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09952_ (.I(_01786_),
    .Z(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09953_ (.A1(\channels.freq3[11] ),
    .A2(_02252_),
    .B(_02255_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09954_ (.A1(_02259_),
    .A2(_02251_),
    .B(_02260_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09955_ (.I(_02250_),
    .Z(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09956_ (.I(_02250_),
    .Z(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09957_ (.A1(\channels.freq3[12] ),
    .A2(_02262_),
    .B(_02255_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09958_ (.A1(_02238_),
    .A2(_02261_),
    .B(_02263_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09959_ (.I(_01071_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09960_ (.I(_02264_),
    .Z(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09961_ (.I(_02265_),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09962_ (.A1(\channels.freq3[13] ),
    .A2(_02262_),
    .B(_02266_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09963_ (.A1(_02242_),
    .A2(_02261_),
    .B(_02267_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09964_ (.A1(\channels.freq3[14] ),
    .A2(_02262_),
    .B(_02266_),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09965_ (.A1(_02245_),
    .A2(_02261_),
    .B(_02268_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09966_ (.A1(\channels.freq3[15] ),
    .A2(_02262_),
    .B(_02266_),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09967_ (.A1(_02247_),
    .A2(_02261_),
    .B(_02269_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09968_ (.A1(_02100_),
    .A2(_01853_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09969_ (.I(_02270_),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09970_ (.I(_02270_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09971_ (.A1(\channels.pw3[8] ),
    .A2(_02272_),
    .B(_02266_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09972_ (.A1(_02249_),
    .A2(_02271_),
    .B(_02273_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09973_ (.I(_02265_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09974_ (.A1(\channels.pw3[9] ),
    .A2(_02272_),
    .B(_02274_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09975_ (.A1(_02254_),
    .A2(_02271_),
    .B(_02275_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09976_ (.A1(\channels.pw3[10] ),
    .A2(_02272_),
    .B(_02274_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09977_ (.A1(_02257_),
    .A2(_02271_),
    .B(_02276_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09978_ (.A1(\channels.pw3[11] ),
    .A2(_02272_),
    .B(_02274_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09979_ (.A1(_02259_),
    .A2(_02271_),
    .B(_02277_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09980_ (.A1(_02229_),
    .A2(_01891_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09981_ (.I(_02278_),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09982_ (.I(_02278_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09983_ (.A1(\channels.ctrl_reg3[0] ),
    .A2(_02280_),
    .B(_02274_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09984_ (.A1(_02249_),
    .A2(_02279_),
    .B(_02281_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09985_ (.I(_02265_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09986_ (.A1(\channels.ctrl_reg3[1] ),
    .A2(_02280_),
    .B(_02282_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09987_ (.A1(_02254_),
    .A2(_02279_),
    .B(_02283_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09988_ (.A1(\channels.ctrl_reg3[2] ),
    .A2(_02280_),
    .B(_02282_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09989_ (.A1(_02257_),
    .A2(_02279_),
    .B(_02284_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09990_ (.A1(\channels.ctrl_reg3[3] ),
    .A2(_02280_),
    .B(_02282_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09991_ (.A1(_02259_),
    .A2(_02279_),
    .B(_02285_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09992_ (.I(_02278_),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09993_ (.I(_02278_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09994_ (.A1(\channels.ctrl_reg3[4] ),
    .A2(_02287_),
    .B(_02282_),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09995_ (.A1(_02238_),
    .A2(_02286_),
    .B(_02288_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09996_ (.I(_02265_),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09997_ (.A1(\channels.ctrl_reg3[5] ),
    .A2(_02287_),
    .B(_02289_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09998_ (.A1(_02242_),
    .A2(_02286_),
    .B(_02290_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09999_ (.A1(\channels.ctrl_reg3[6] ),
    .A2(_02287_),
    .B(_02289_),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10000_ (.A1(_02245_),
    .A2(_02286_),
    .B(_02291_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10001_ (.A1(\channels.ctrl_reg3[7] ),
    .A2(_02287_),
    .B(_02289_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10002_ (.A1(_02247_),
    .A2(_02286_),
    .B(_02292_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10003_ (.A1(_02229_),
    .A2(_01876_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10004_ (.I(_02293_),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10005_ (.I(_02293_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10006_ (.A1(\channels.atk_dec3[0] ),
    .A2(_02295_),
    .B(_02289_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10007_ (.A1(_02249_),
    .A2(_02294_),
    .B(_02296_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10008_ (.I(_02264_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10009_ (.I(_02297_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10010_ (.A1(\channels.atk_dec3[1] ),
    .A2(_02295_),
    .B(_02298_),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10011_ (.A1(_02254_),
    .A2(_02294_),
    .B(_02299_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10012_ (.A1(\channels.atk_dec3[2] ),
    .A2(_02295_),
    .B(_02298_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10013_ (.A1(_02257_),
    .A2(_02294_),
    .B(_02300_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10014_ (.A1(\channels.atk_dec3[3] ),
    .A2(_02295_),
    .B(_02298_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10015_ (.A1(_02259_),
    .A2(_02294_),
    .B(_02301_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10016_ (.I(_02293_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10017_ (.I(_02293_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10018_ (.A1(\channels.atk_dec3[4] ),
    .A2(_02303_),
    .B(_02298_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10019_ (.A1(_02238_),
    .A2(_02302_),
    .B(_02304_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10020_ (.I(_02297_),
    .Z(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10021_ (.A1(\channels.atk_dec3[5] ),
    .A2(_02303_),
    .B(_02305_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10022_ (.A1(_02242_),
    .A2(_02302_),
    .B(_02306_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10023_ (.A1(\channels.atk_dec3[6] ),
    .A2(_02303_),
    .B(_02305_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10024_ (.A1(_02245_),
    .A2(_02302_),
    .B(_02307_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10025_ (.A1(\channels.atk_dec3[7] ),
    .A2(_02303_),
    .B(_02305_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10026_ (.A1(_02247_),
    .A2(_02302_),
    .B(_02308_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10027_ (.I(_02109_),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10028_ (.I(_01789_),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10029_ (.A1(_02310_),
    .A2(_01955_),
    .Z(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10030_ (.I(_02311_),
    .Z(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10031_ (.I(_02311_),
    .Z(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10032_ (.A1(\channels.sus_rel3[0] ),
    .A2(_02313_),
    .B(_02305_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10033_ (.A1(_02309_),
    .A2(_02312_),
    .B(_02314_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10034_ (.I(_02188_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10035_ (.I(_02297_),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10036_ (.A1(\channels.sus_rel3[1] ),
    .A2(_02313_),
    .B(_02316_),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10037_ (.A1(_02315_),
    .A2(_02312_),
    .B(_02317_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10038_ (.I(_02193_),
    .Z(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10039_ (.A1(\channels.sus_rel3[2] ),
    .A2(_02313_),
    .B(_02316_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10040_ (.A1(_02318_),
    .A2(_02312_),
    .B(_02319_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10041_ (.I(_01785_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10042_ (.I(_02320_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10043_ (.A1(\channels.sus_rel3[3] ),
    .A2(_02313_),
    .B(_02316_),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10044_ (.A1(_02321_),
    .A2(_02312_),
    .B(_02322_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10045_ (.I(_02311_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10046_ (.I(_02311_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10047_ (.A1(\channels.sus_rel3[4] ),
    .A2(_02324_),
    .B(_02316_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10048_ (.A1(_01805_),
    .A2(_02323_),
    .B(_02325_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10049_ (.I(_02160_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10050_ (.I(_02297_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10051_ (.A1(\channels.sus_rel3[5] ),
    .A2(_02324_),
    .B(_02327_),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10052_ (.A1(_02326_),
    .A2(_02323_),
    .B(_02328_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10053_ (.I(_01817_),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10054_ (.A1(\channels.sus_rel3[6] ),
    .A2(_02324_),
    .B(_02327_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10055_ (.A1(_02329_),
    .A2(_02323_),
    .B(_02330_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10056_ (.I(_01822_),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10057_ (.A1(\channels.sus_rel3[7] ),
    .A2(_02324_),
    .B(_02327_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10058_ (.A1(_02331_),
    .A2(_02323_),
    .B(_02332_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10059_ (.A1(_02310_),
    .A2(_01968_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10060_ (.I(_02333_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10061_ (.I(_02333_),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10062_ (.A1(\filters.cutoff_lut[9] ),
    .A2(_02335_),
    .B(_02327_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10063_ (.A1(_02309_),
    .A2(_02334_),
    .B(_02336_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10064_ (.I(_02264_),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10065_ (.I(_02337_),
    .Z(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10066_ (.A1(\filters.cutoff_lut[10] ),
    .A2(_02335_),
    .B(_02338_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10067_ (.A1(_02315_),
    .A2(_02334_),
    .B(_02339_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10068_ (.A1(\filters.cutoff_lut[11] ),
    .A2(_02335_),
    .B(_02338_),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10069_ (.A1(_02318_),
    .A2(_02334_),
    .B(_02340_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10070_ (.A1(\filters.cutoff_lut[12] ),
    .A2(_02335_),
    .B(_02338_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10071_ (.A1(_02321_),
    .A2(_02334_),
    .B(_02341_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10072_ (.I(_02333_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10073_ (.I(_02333_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10074_ (.A1(\filters.cutoff_lut[13] ),
    .A2(_02343_),
    .B(_02338_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10075_ (.A1(_01805_),
    .A2(_02342_),
    .B(_02344_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10076_ (.I(_02337_),
    .Z(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10077_ (.A1(\filters.cutoff_lut[14] ),
    .A2(_02343_),
    .B(_02345_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10078_ (.A1(_02326_),
    .A2(_02342_),
    .B(_02346_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10079_ (.A1(\filters.cutoff_lut[15] ),
    .A2(_02343_),
    .B(_02345_),
    .ZN(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10080_ (.A1(_02329_),
    .A2(_02342_),
    .B(_02347_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10081_ (.A1(\filters.cutoff_lut[16] ),
    .A2(_02343_),
    .B(_02345_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10082_ (.A1(_02331_),
    .A2(_02342_),
    .B(_02348_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10083_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.in ),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _10084_ (.I0(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ),
    .I1(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ),
    .I2(\tt_um_rejunity_sn76489.noise[0].gen.counter[6] ),
    .I3(_02349_),
    .S0(\tt_um_rejunity_sn76489.control_noise[0][0] ),
    .S1(\tt_um_rejunity_sn76489.control_noise[0][1] ),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10085_ (.I(_02350_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10086_ (.A1(_01945_),
    .A2(_02351_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10087_ (.I(_01790_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10088_ (.A1(_02352_),
    .A2(_01917_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10089_ (.A1(net7),
    .A2(_02353_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10090_ (.I(_01826_),
    .Z(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10091_ (.I(_02355_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10092_ (.A1(_01075_),
    .A2(_02353_),
    .B(_02354_),
    .C(_02356_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10093_ (.A1(net8),
    .A2(_02353_),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10094_ (.A1(_01076_),
    .A2(_02353_),
    .B(_02357_),
    .C(_02356_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10095_ (.I(_01093_),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10096_ (.A1(_01081_),
    .A2(_02358_),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10097_ (.I(_02359_),
    .Z(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10098_ (.I(_02360_),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10099_ (.I(_01096_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10100_ (.A1(_02362_),
    .A2(_01579_),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10101_ (.A1(\channels.sync_outs[2] ),
    .A2(_01255_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10102_ (.A1(_02361_),
    .A2(_02363_),
    .B(_02364_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10103_ (.I(_01292_),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10104_ (.A1(_01081_),
    .A2(_02365_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10105_ (.I(_02366_),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10106_ (.I(_02367_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10107_ (.A1(\channels.sync_outs[1] ),
    .A2(_01240_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10108_ (.A1(_02368_),
    .A2(_02363_),
    .B(_02369_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10109_ (.A1(\channels.sync_outs[0] ),
    .A2(_01570_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10110_ (.A1(_01550_),
    .A2(_02363_),
    .B(_02370_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10111_ (.A1(_01277_),
    .A2(\channels.ctrl_reg2[4] ),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10112_ (.A1(_01276_),
    .A2(\channels.ctrl_reg3[4] ),
    .B1(\channels.ctrl_reg1[4] ),
    .B2(_01262_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10113_ (.A1(_01274_),
    .A2(_02371_),
    .B(_02372_),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10114_ (.I(_02373_),
    .Z(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10115_ (.A1(\channels.ctrl_reg2[2] ),
    .A2(\channels.ring_outs[0] ),
    .A3(_01283_),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10116_ (.A1(\channels.ctrl_reg3[2] ),
    .A2(\channels.ring_outs[1] ),
    .A3(_01084_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10117_ (.A1(\channels.ctrl_reg1[2] ),
    .A2(\channels.ring_outs[2] ),
    .A3(_01294_),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10118_ (.A1(_02375_),
    .A2(_02376_),
    .A3(_02377_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10119_ (.A1(_02362_),
    .A2(_02378_),
    .Z(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10120_ (.I(_02379_),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10121_ (.A1(_01537_),
    .A2(_02380_),
    .Z(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10122_ (.A1(\channels.ctrl_reg1[5] ),
    .A2(_01296_),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10123_ (.A1(\channels.ctrl_reg3[5] ),
    .A2(_01085_),
    .B1(_01284_),
    .B2(\channels.ctrl_reg2[5] ),
    .C(_02382_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10124_ (.I(_02383_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10125_ (.A1(\channels.ctrl_reg3[7] ),
    .A2(_01084_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10126_ (.A1(\channels.ctrl_reg2[7] ),
    .A2(_01283_),
    .B1(_01296_),
    .B2(\channels.ctrl_reg1[7] ),
    .ZN(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10127_ (.A1(_02385_),
    .A2(_02386_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10128_ (.I(_02387_),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10129_ (.A1(_01643_),
    .A2(_02388_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10130_ (.A1(_01544_),
    .A2(_02384_),
    .B(_02389_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10131_ (.I(_01258_),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10132_ (.I(_01282_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10133_ (.A1(_02391_),
    .A2(_02392_),
    .A3(\channels.pw3[11] ),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10134_ (.A1(_02392_),
    .A2(\channels.pw2[11] ),
    .B(_01107_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10135_ (.A1(\channels.pw1[11] ),
    .A2(_01261_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10136_ (.A1(_02393_),
    .A2(_02394_),
    .B(_02395_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10137_ (.A1(_02362_),
    .A2(_02396_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10138_ (.A1(_02393_),
    .A2(_02394_),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10139_ (.I(_01082_),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10140_ (.A1(_02399_),
    .A2(_01260_),
    .A3(\channels.pw2[10] ),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10141_ (.A1(_02391_),
    .A2(_02392_),
    .A3(\channels.pw3[10] ),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10142_ (.A1(\channels.pw1[10] ),
    .A2(_01295_),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10143_ (.A1(_02400_),
    .A2(_02401_),
    .A3(_02402_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _10144_ (.I0(\channels.accum[0][22] ),
    .I1(\channels.accum[1][22] ),
    .I2(\channels.accum[2][22] ),
    .I3(\channels.accum[3][22] ),
    .S0(_01505_),
    .S1(_01506_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _10145_ (.A1(_01096_),
    .A2(_02398_),
    .A3(_02395_),
    .B1(_02403_),
    .B2(_02404_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10146_ (.I(_01565_),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10147_ (.I(_01282_),
    .Z(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10148_ (.A1(_02391_),
    .A2(_02407_),
    .A3(\channels.pw3[9] ),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10149_ (.A1(_02392_),
    .A2(\channels.pw2[9] ),
    .B(_02399_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10150_ (.A1(\channels.pw1[9] ),
    .A2(_01261_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10151_ (.A1(_02408_),
    .A2(_02409_),
    .B(_02410_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10152_ (.A1(_02399_),
    .A2(_01260_),
    .A3(\channels.pw2[8] ),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10153_ (.A1(_02391_),
    .A2(_02407_),
    .A3(\channels.pw3[8] ),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10154_ (.A1(\channels.pw1[8] ),
    .A2(_01295_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10155_ (.A1(_02412_),
    .A2(_02413_),
    .A3(_02414_),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10156_ (.A1(_02406_),
    .A2(_02411_),
    .B1(_02415_),
    .B2(_01563_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10157_ (.A1(_02400_),
    .A2(_02401_),
    .A3(_02402_),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10158_ (.A1(_01576_),
    .A2(_02417_),
    .B1(_02411_),
    .B2(_02406_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10159_ (.A1(_02416_),
    .A2(_02418_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10160_ (.A1(_02405_),
    .A2(_02419_),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10161_ (.A1(_02408_),
    .A2(_02409_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10162_ (.A1(_02412_),
    .A2(_02413_),
    .A3(_02414_),
    .Z(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10163_ (.A1(_01565_),
    .A2(_02421_),
    .A3(_02410_),
    .B1(_02422_),
    .B2(_01560_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10164_ (.A1(_02362_),
    .A2(_02396_),
    .B1(_02415_),
    .B2(_01563_),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10165_ (.A1(_02405_),
    .A2(_02423_),
    .A3(_02418_),
    .A4(_02424_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10166_ (.I(_02425_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10167_ (.A1(_01108_),
    .A2(_01109_),
    .A3(\channels.pw2[7] ),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10168_ (.I(_01259_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10169_ (.I(_01282_),
    .Z(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10170_ (.I(_02429_),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10171_ (.A1(_02428_),
    .A2(_02430_),
    .A3(\channels.pw3[7] ),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10172_ (.I(_01294_),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10173_ (.A1(\channels.pw1[7] ),
    .A2(_02432_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10174_ (.A1(_01551_),
    .A2(_02427_),
    .A3(_02431_),
    .A4(_02433_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _10175_ (.A1(_02427_),
    .A2(_02431_),
    .A3(_02433_),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10176_ (.I(\channels.pw1[5] ),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10177_ (.I(_01295_),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10178_ (.A1(_02428_),
    .A2(_02407_),
    .A3(\channels.pw3[5] ),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10179_ (.A1(_02430_),
    .A2(\channels.pw2[5] ),
    .B(_01108_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10180_ (.A1(_02436_),
    .A2(_02437_),
    .B1(_02438_),
    .B2(_02439_),
    .C(_01537_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10181_ (.I(\channels.pw1[4] ),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10182_ (.A1(_02428_),
    .A2(_02430_),
    .A3(\channels.pw3[4] ),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10183_ (.A1(_02430_),
    .A2(\channels.pw2[4] ),
    .B(_01108_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10184_ (.A1(_02441_),
    .A2(_01296_),
    .B1(_02442_),
    .B2(_02443_),
    .C(_01530_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10185_ (.A1(_02440_),
    .A2(_02444_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10186_ (.A1(_02399_),
    .A2(_01109_),
    .A3(\channels.pw2[6] ),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10187_ (.A1(_02428_),
    .A2(_02407_),
    .A3(\channels.pw3[6] ),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10188_ (.A1(\channels.pw1[6] ),
    .A2(_02432_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10189_ (.A1(_01543_),
    .A2(_02446_),
    .A3(_02447_),
    .A4(_02448_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10190_ (.A1(_01275_),
    .A2(_01273_),
    .A3(\channels.pw2[5] ),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10191_ (.A1(\channels.pw1[5] ),
    .A2(_02437_),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10192_ (.A1(_01537_),
    .A2(_02450_),
    .A3(_02438_),
    .A4(_02451_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _10193_ (.A1(_02449_),
    .A2(_02452_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _10194_ (.A1(_02446_),
    .A2(_02447_),
    .A3(_02448_),
    .Z(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _10195_ (.A1(_01551_),
    .A2(_02435_),
    .B1(_02445_),
    .B2(_02453_),
    .C1(_02454_),
    .C2(_01543_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10196_ (.I(\channels.pw2[2] ),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10197_ (.I(_02429_),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10198_ (.A1(_01592_),
    .A2(_02457_),
    .A3(\channels.pw3[2] ),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10199_ (.A1(\channels.pw1[2] ),
    .A2(_02432_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10200_ (.A1(_02456_),
    .A2(_01110_),
    .B(_02458_),
    .C(_02459_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10201_ (.A1(_01508_),
    .A2(_02460_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10202_ (.A1(_01275_),
    .A2(_01273_),
    .A3(\channels.pw2[0] ),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10203_ (.A1(_01592_),
    .A2(_02457_),
    .A3(\channels.pw3[0] ),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10204_ (.A1(\channels.pw1[0] ),
    .A2(_02437_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10205_ (.A1(_01479_),
    .A2(_02462_),
    .A3(_02463_),
    .A4(_02464_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10206_ (.A1(_01259_),
    .A2(_02429_),
    .A3(\channels.pw3[1] ),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10207_ (.A1(_01083_),
    .A2(\channels.pw1[1] ),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10208_ (.A1(_02429_),
    .A2(\channels.pw2[1] ),
    .B(_02467_),
    .C(_01107_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10209_ (.A1(_01491_),
    .A2(_02466_),
    .A3(_02468_),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10210_ (.A1(_02466_),
    .A2(_02468_),
    .B(_01491_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10211_ (.A1(_02465_),
    .A2(_02469_),
    .B(_02470_),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10212_ (.I(\channels.pw2[3] ),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10213_ (.A1(_01592_),
    .A2(_02457_),
    .A3(\channels.pw3[3] ),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10214_ (.A1(\channels.pw1[3] ),
    .A2(_02432_),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10215_ (.A1(_02472_),
    .A2(_01110_),
    .B(_02473_),
    .C(_02474_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10216_ (.A1(_01519_),
    .A2(_02475_),
    .B1(_02460_),
    .B2(_01508_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10217_ (.A1(_02461_),
    .A2(_02471_),
    .B(_02476_),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _10218_ (.A1(_01551_),
    .A2(_02435_),
    .B1(_02454_),
    .B2(_01543_),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _10219_ (.A1(_02440_),
    .A2(_02444_),
    .Z(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10220_ (.A1(_01275_),
    .A2(_01109_),
    .A3(\channels.pw2[4] ),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10221_ (.A1(\channels.pw1[4] ),
    .A2(_02437_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10222_ (.A1(_01530_),
    .A2(_02480_),
    .A3(_02442_),
    .A4(_02481_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10223_ (.A1(_01519_),
    .A2(_02475_),
    .B(_02482_),
    .C(_02434_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10224_ (.A1(_02478_),
    .A2(_02479_),
    .A3(_02453_),
    .A4(_02483_),
    .ZN(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10225_ (.A1(_02434_),
    .A2(_02455_),
    .B1(_02477_),
    .B2(_02484_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _10226_ (.A1(_02397_),
    .A2(_02420_),
    .B1(_02426_),
    .B2(_02485_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10227_ (.A1(_02434_),
    .A2(_02482_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10228_ (.A1(_02478_),
    .A2(_02479_),
    .A3(_02453_),
    .A4(_02487_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10229_ (.A1(_02466_),
    .A2(_02468_),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10230_ (.A1(_01491_),
    .A2(_02489_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10231_ (.A1(_02465_),
    .A2(_02490_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10232_ (.A1(_01520_),
    .A2(_02475_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10233_ (.A1(_02463_),
    .A2(_02464_),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10234_ (.A1(_02462_),
    .A2(_02493_),
    .B(_01479_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10235_ (.A1(_02461_),
    .A2(_02492_),
    .A3(_02494_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10236_ (.A1(_02425_),
    .A2(_02476_),
    .A3(_02491_),
    .A4(_02495_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10237_ (.A1(_01276_),
    .A2(\channels.ctrl_reg2[6] ),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10238_ (.A1(_01273_),
    .A2(_02497_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _10239_ (.A1(_01276_),
    .A2(\channels.ctrl_reg3[6] ),
    .B1(\channels.ctrl_reg1[6] ),
    .B2(_01262_),
    .C(_02498_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10240_ (.A1(_02488_),
    .A2(_02496_),
    .B(_02499_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10241_ (.A1(_02486_),
    .A2(_02500_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10242_ (.A1(_02374_),
    .A2(_02381_),
    .B(_02390_),
    .C(_02501_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10243_ (.I(_02502_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10244_ (.I(_02503_),
    .Z(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _10245_ (.I0(\channels.env_vol[0][0] ),
    .I1(\channels.env_vol[1][0] ),
    .I2(\channels.ch3_env[0] ),
    .I3(\channels.env_vol[3][0] ),
    .S0(_01155_),
    .S1(_01169_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10246_ (.I(_02505_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10247_ (.I(_02506_),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10248_ (.A1(_02504_),
    .A2(_02507_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10249_ (.A1(_02486_),
    .A2(_02500_),
    .B(_02388_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10250_ (.I(_02509_),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10251_ (.I(_02510_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10252_ (.A1(_01507_),
    .A2(_02380_),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10253_ (.A1(_01518_),
    .A2(_02383_),
    .ZN(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10254_ (.A1(_02374_),
    .A2(_02512_),
    .B(_02513_),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10255_ (.I(_02514_),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10256_ (.I(_02515_),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10257_ (.I(\channels.ch3_env[2] ),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10258_ (.A1(_01316_),
    .A2(_02517_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10259_ (.A1(_01316_),
    .A2(\channels.env_vol[3][2] ),
    .B(_02518_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10260_ (.I(_01151_),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10261_ (.I(_02520_),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10262_ (.I0(\channels.env_vol[0][2] ),
    .I1(\channels.env_vol[1][2] ),
    .S(_02521_),
    .Z(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10263_ (.A1(_01167_),
    .A2(_02522_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10264_ (.A1(_01699_),
    .A2(_02519_),
    .B(_02523_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10265_ (.A1(_02511_),
    .A2(_02516_),
    .A3(_02524_),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10266_ (.I(_02510_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10267_ (.A1(_01492_),
    .A2(_02380_),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10268_ (.A1(_01507_),
    .A2(_02384_),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10269_ (.A1(_02374_),
    .A2(_02527_),
    .B(_02528_),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10270_ (.I(_02529_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10271_ (.I(_01667_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10272_ (.I(\channels.ch3_env[3] ),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10273_ (.A1(_01315_),
    .A2(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10274_ (.A1(_01153_),
    .A2(\channels.env_vol[3][3] ),
    .B(_02533_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10275_ (.I0(\channels.env_vol[0][3] ),
    .I1(\channels.env_vol[1][3] ),
    .S(_02520_),
    .Z(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10276_ (.A1(_01166_),
    .A2(_02535_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10277_ (.A1(_02531_),
    .A2(_02534_),
    .B(_02536_),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10278_ (.I(_02537_),
    .Z(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10279_ (.A1(_02526_),
    .A2(_02530_),
    .A3(_02538_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10280_ (.I(_02374_),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10281_ (.I(_02380_),
    .Z(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10282_ (.A1(_01480_),
    .A2(_02541_),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10283_ (.I(_02384_),
    .Z(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10284_ (.A1(_01492_),
    .A2(_02543_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10285_ (.A1(_02540_),
    .A2(_02542_),
    .B(_02544_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _10286_ (.I0(\channels.env_vol[0][4] ),
    .I1(\channels.env_vol[1][4] ),
    .I2(\channels.ch3_env[4] ),
    .I3(\channels.env_vol[3][4] ),
    .S0(_01153_),
    .S1(_01698_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10287_ (.A1(_02526_),
    .A2(_02545_),
    .A3(_02546_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10288_ (.A1(_02539_),
    .A2(_02547_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10289_ (.A1(_02539_),
    .A2(_02547_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10290_ (.A1(_02525_),
    .A2(_02548_),
    .B(_02549_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10291_ (.A1(_01531_),
    .A2(_02379_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10292_ (.I(_02373_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10293_ (.A1(_01626_),
    .A2(_02387_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10294_ (.A1(_01538_),
    .A2(_02384_),
    .B1(_02551_),
    .B2(_02552_),
    .C(_02553_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10295_ (.A1(_02486_),
    .A2(_02500_),
    .B(_02554_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10296_ (.I(_02555_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10297_ (.I(_02556_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10298_ (.I(\channels.ch3_env[1] ),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10299_ (.A1(_01317_),
    .A2(_02558_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10300_ (.A1(_01317_),
    .A2(\channels.env_vol[3][1] ),
    .B(_02559_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10301_ (.I0(\channels.env_vol[0][1] ),
    .I1(\channels.env_vol[1][1] ),
    .S(_01154_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10302_ (.A1(_01338_),
    .A2(_02561_),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10303_ (.A1(_01338_),
    .A2(_02560_),
    .B(_02562_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10304_ (.I(_02563_),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10305_ (.A1(_02557_),
    .A2(_02564_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10306_ (.A1(_02550_),
    .A2(_02565_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10307_ (.A1(_02550_),
    .A2(_02565_),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10308_ (.A1(_02508_),
    .A2(_02566_),
    .B(_02567_),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10309_ (.I(_02541_),
    .Z(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10310_ (.A1(_01480_),
    .A2(_02543_),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10311_ (.A1(_02569_),
    .A2(_02540_),
    .B(_02570_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10312_ (.I(\channels.ch3_env[6] ),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10313_ (.A1(_02520_),
    .A2(_02572_),
    .ZN(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10314_ (.A1(_02521_),
    .A2(\channels.env_vol[3][6] ),
    .B(_02573_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10315_ (.I0(\channels.env_vol[0][6] ),
    .I1(\channels.env_vol[1][6] ),
    .S(_01152_),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10316_ (.A1(_01166_),
    .A2(_02575_),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10317_ (.A1(_01698_),
    .A2(_02574_),
    .B(_02576_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10318_ (.I(_02577_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10319_ (.A1(_02526_),
    .A2(_02571_),
    .A3(_02578_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10320_ (.I(\channels.ch3_env[5] ),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10321_ (.A1(_01153_),
    .A2(_02580_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10322_ (.A1(_01316_),
    .A2(\channels.env_vol[3][5] ),
    .B(_02581_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10323_ (.I0(\channels.env_vol[0][5] ),
    .I1(\channels.env_vol[1][5] ),
    .S(_02521_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10324_ (.A1(_01167_),
    .A2(_02583_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10325_ (.A1(_01699_),
    .A2(_02582_),
    .B(_02584_),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10326_ (.A1(_02526_),
    .A2(_02545_),
    .A3(_02585_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10327_ (.A1(_02579_),
    .A2(_02586_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10328_ (.A1(_01520_),
    .A2(_02379_),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10329_ (.A1(_01609_),
    .A2(_02387_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10330_ (.A1(_01531_),
    .A2(_02383_),
    .B1(_02588_),
    .B2(_02552_),
    .C(_02589_),
    .ZN(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10331_ (.A1(_02486_),
    .A2(_02500_),
    .B(_02590_),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10332_ (.I(_02591_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10333_ (.A1(_02524_),
    .A2(_02592_),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10334_ (.I(_02509_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10335_ (.A1(_02594_),
    .A2(_02537_),
    .A3(_02515_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10336_ (.I(_02546_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10337_ (.A1(_02511_),
    .A2(_02530_),
    .A3(_02596_),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10338_ (.A1(_02593_),
    .A2(_02595_),
    .A3(_02597_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10339_ (.A1(_02587_),
    .A2(_02598_),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10340_ (.I(_02594_),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10341_ (.I(_02600_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10342_ (.I(_02571_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10343_ (.I(_02585_),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10344_ (.I(_02603_),
    .Z(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10345_ (.A1(_02601_),
    .A2(_02602_),
    .A3(_02604_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10346_ (.A1(_02539_),
    .A2(_02547_),
    .A3(_02525_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10347_ (.A1(_02605_),
    .A2(_02606_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10348_ (.A1(_02599_),
    .A2(_02607_),
    .ZN(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10349_ (.I(_02505_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10350_ (.A1(_02504_),
    .A2(_02609_),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10351_ (.A1(_02550_),
    .A2(_02565_),
    .A3(_02610_),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10352_ (.A1(_02599_),
    .A2(_02607_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10353_ (.A1(_02608_),
    .A2(_02611_),
    .B(_02612_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10354_ (.A1(_02587_),
    .A2(_02598_),
    .ZN(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10355_ (.I(_02593_),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10356_ (.A1(_02595_),
    .A2(_02597_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10357_ (.A1(_02595_),
    .A2(_02597_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10358_ (.A1(_02615_),
    .A2(_02616_),
    .B(_02617_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10359_ (.A1(_02564_),
    .A2(_02504_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10360_ (.A1(_02618_),
    .A2(_02619_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10361_ (.A1(_01544_),
    .A2(_02541_),
    .Z(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10362_ (.A1(_01668_),
    .A2(_02388_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10363_ (.A1(_01552_),
    .A2(_02543_),
    .B(_02622_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10364_ (.A1(_02540_),
    .A2(_02621_),
    .B(_02623_),
    .C(_02501_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10365_ (.I(_02624_),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10366_ (.I(_02625_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10367_ (.A1(_02506_),
    .A2(_02626_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10368_ (.A1(_02620_),
    .A2(_02627_),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10369_ (.A1(_02579_),
    .A2(_02586_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10370_ (.I(_02530_),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10371_ (.A1(_02600_),
    .A2(_02630_),
    .A3(_02603_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10372_ (.I(_02545_),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10373_ (.A1(_02600_),
    .A2(_02632_),
    .A3(_02578_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10374_ (.I(\channels.ch3_env[7] ),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10375_ (.A1(_01315_),
    .A2(_02634_),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10376_ (.A1(_02521_),
    .A2(\channels.env_vol[3][7] ),
    .B(_02635_),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10377_ (.I0(\channels.env_vol[0][7] ),
    .I1(\channels.env_vol[1][7] ),
    .S(_02520_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10378_ (.A1(_01166_),
    .A2(_02637_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10379_ (.A1(_02531_),
    .A2(_02636_),
    .B(_02638_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10380_ (.I(_02639_),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10381_ (.A1(_02511_),
    .A2(_02571_),
    .A3(_02640_),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10382_ (.A1(_02631_),
    .A2(_02633_),
    .A3(_02641_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10383_ (.I(_02524_),
    .Z(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10384_ (.I(_02643_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10385_ (.A1(_02644_),
    .A2(_02557_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10386_ (.I(_02538_),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10387_ (.I(_02592_),
    .Z(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10388_ (.A1(_02646_),
    .A2(_02647_),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10389_ (.A1(_02511_),
    .A2(_02596_),
    .A3(_02515_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10390_ (.A1(_02648_),
    .A2(_02649_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10391_ (.A1(_02645_),
    .A2(_02650_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10392_ (.A1(_02629_),
    .A2(_02642_),
    .A3(_02651_),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10393_ (.A1(_02614_),
    .A2(_02628_),
    .A3(_02652_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10394_ (.A1(_02568_),
    .A2(_02613_),
    .A3(_02653_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10395_ (.A1(_02557_),
    .A2(_02505_),
    .Z(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10396_ (.A1(_02601_),
    .A2(_02630_),
    .A3(_02644_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10397_ (.I(_02600_),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10398_ (.A1(_02657_),
    .A2(_02646_),
    .A3(_02632_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10399_ (.I(_02546_),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10400_ (.A1(_02657_),
    .A2(_02659_),
    .A3(_02571_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10401_ (.A1(_02658_),
    .A2(_02660_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10402_ (.A1(_02658_),
    .A2(_02660_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10403_ (.A1(_02656_),
    .A2(_02661_),
    .B(_02662_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10404_ (.I(_02563_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10405_ (.A1(_02664_),
    .A2(_02647_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10406_ (.A1(_02663_),
    .A2(_02665_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10407_ (.A1(_02663_),
    .A2(_02665_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10408_ (.A1(_02655_),
    .A2(_02666_),
    .B(_02667_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10409_ (.A1(_02605_),
    .A2(_02606_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10410_ (.A1(_02655_),
    .A2(_02663_),
    .A3(_02665_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10411_ (.A1(_02669_),
    .A2(_02670_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10412_ (.A1(_02608_),
    .A2(_02611_),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10413_ (.A1(_02671_),
    .A2(_02672_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10414_ (.A1(_02671_),
    .A2(_02672_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10415_ (.A1(_02668_),
    .A2(_02673_),
    .B(_02674_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10416_ (.A1(_02669_),
    .A2(_02670_),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10417_ (.A1(_02601_),
    .A2(_02516_),
    .A3(_02664_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10418_ (.I(_02646_),
    .Z(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10419_ (.A1(_02657_),
    .A2(_02678_),
    .A3(_02602_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10420_ (.A1(_02657_),
    .A2(_02632_),
    .A3(_02643_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10421_ (.A1(_02679_),
    .A2(_02680_),
    .ZN(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10422_ (.A1(_02609_),
    .A2(_02647_),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _10423_ (.A1(_02677_),
    .A2(_02681_),
    .A3(_02682_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _10424_ (.A1(_02658_),
    .A2(_02660_),
    .A3(_02656_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10425_ (.A1(_02671_),
    .A2(_02676_),
    .A3(_02683_),
    .A4(_02684_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10426_ (.I(_02601_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10427_ (.I(_02686_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10428_ (.I(_02564_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10429_ (.I(_02688_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10430_ (.A1(_02687_),
    .A2(_02516_),
    .A3(_02689_),
    .A4(_02681_),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10431_ (.A1(_02677_),
    .A2(_02681_),
    .Z(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10432_ (.A1(_02691_),
    .A2(_02682_),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10433_ (.A1(_02683_),
    .A2(_02684_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10434_ (.A1(_02669_),
    .A2(_02670_),
    .A3(_02693_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10435_ (.A1(_02690_),
    .A2(_02692_),
    .B(_02694_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10436_ (.A1(_02671_),
    .A2(_02672_),
    .A3(_02668_),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10437_ (.A1(_02685_),
    .A2(_02695_),
    .B(_02696_),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10438_ (.A1(_02683_),
    .A2(_02684_),
    .Z(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10439_ (.A1(_02686_),
    .A2(_02630_),
    .A3(_02688_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10440_ (.A1(_02686_),
    .A2(_02516_),
    .A3(_02609_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10441_ (.A1(_02699_),
    .A2(_02700_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10442_ (.A1(_02679_),
    .A2(_02680_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10443_ (.A1(_02699_),
    .A2(_02700_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10444_ (.A1(_02701_),
    .A2(_02702_),
    .B(_02703_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10445_ (.I(_02507_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10446_ (.A1(_02686_),
    .A2(_02632_),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10447_ (.A1(_01172_),
    .A2(_02560_),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10448_ (.A1(_01172_),
    .A2(_02561_),
    .B(_02707_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10449_ (.I(_02708_),
    .Z(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10450_ (.A1(_02706_),
    .A2(_02709_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10451_ (.A1(_02687_),
    .A2(_02630_),
    .A3(_02705_),
    .A4(_02710_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10452_ (.I(_02644_),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _10453_ (.I(_02507_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10454_ (.A1(_02510_),
    .A2(_02529_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10455_ (.I(_02714_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10456_ (.A1(_02706_),
    .A2(_02708_),
    .B1(_02713_),
    .B2(_02715_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10457_ (.A1(_02687_),
    .A2(_02712_),
    .A3(_02602_),
    .A4(_02716_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10458_ (.A1(_02701_),
    .A2(_02702_),
    .ZN(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10459_ (.A1(_02711_),
    .A2(_02717_),
    .B(_02718_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10460_ (.A1(_02683_),
    .A2(_02684_),
    .A3(_02704_),
    .Z(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10461_ (.A1(_02719_),
    .A2(_02720_),
    .Z(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10462_ (.A1(_01174_),
    .A2(_02519_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10463_ (.A1(_01174_),
    .A2(_02522_),
    .B(_02722_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10464_ (.A1(_02715_),
    .A2(_02723_),
    .B(_02718_),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10465_ (.A1(_02687_),
    .A2(_02705_),
    .A3(_02602_),
    .A4(_02710_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10466_ (.A1(_02656_),
    .A2(_02718_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10467_ (.A1(_02719_),
    .A2(_02720_),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10468_ (.A1(_02724_),
    .A2(_02725_),
    .A3(_02726_),
    .B(_02727_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10469_ (.A1(_02698_),
    .A2(_02704_),
    .B1(_02721_),
    .B2(_02728_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10470_ (.A1(_02690_),
    .A2(_02692_),
    .A3(_02694_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10471_ (.A1(_02685_),
    .A2(_02695_),
    .A3(_02696_),
    .B(_02730_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10472_ (.A1(_02695_),
    .A2(_02729_),
    .A3(_02731_),
    .Z(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10473_ (.A1(_02654_),
    .A2(_02675_),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10474_ (.A1(_02697_),
    .A2(_02732_),
    .B(_02733_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10475_ (.A1(_02654_),
    .A2(_02675_),
    .B(_02734_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10476_ (.A1(_02613_),
    .A2(_02653_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10477_ (.A1(_02613_),
    .A2(_02653_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10478_ (.A1(_02568_),
    .A2(_02736_),
    .B(_02737_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10479_ (.A1(_02705_),
    .A2(_02620_),
    .A3(_02626_),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10480_ (.A1(_02618_),
    .A2(_02619_),
    .B(_02739_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10481_ (.A1(_02614_),
    .A2(_02652_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10482_ (.A1(_02614_),
    .A2(_02652_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10483_ (.A1(_02628_),
    .A2(_02741_),
    .B(_02742_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10484_ (.A1(_02629_),
    .A2(_02642_),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10485_ (.A1(_02629_),
    .A2(_02642_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10486_ (.A1(_02744_),
    .A2(_02651_),
    .B(_02745_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10487_ (.A1(_02633_),
    .A2(_02641_),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10488_ (.A1(_02633_),
    .A2(_02641_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10489_ (.A1(_02631_),
    .A2(_02747_),
    .B(_02748_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10490_ (.A1(_02594_),
    .A2(_02545_),
    .A3(_02640_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10491_ (.A1(_02594_),
    .A2(_02530_),
    .A3(_02578_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10492_ (.A1(_02509_),
    .A2(_02514_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10493_ (.A1(_01699_),
    .A2(_02582_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10494_ (.A1(_01168_),
    .A2(_02583_),
    .B(_02753_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10495_ (.A1(_02752_),
    .A2(_02754_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10496_ (.A1(_02750_),
    .A2(_02751_),
    .A3(_02755_),
    .Z(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10497_ (.A1(_02643_),
    .A2(_02503_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10498_ (.A1(_02596_),
    .A2(_02647_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10499_ (.A1(_02538_),
    .A2(_02556_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10500_ (.A1(_02758_),
    .A2(_02759_),
    .Z(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10501_ (.A1(_02758_),
    .A2(_02759_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10502_ (.A1(_02760_),
    .A2(_02761_),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10503_ (.A1(_02757_),
    .A2(_02762_),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10504_ (.A1(_02749_),
    .A2(_02756_),
    .A3(_02763_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10505_ (.A1(_02746_),
    .A2(_02764_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10506_ (.A1(_02648_),
    .A2(_02649_),
    .Z(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10507_ (.A1(_02645_),
    .A2(_02650_),
    .B(_02766_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10508_ (.A1(_02664_),
    .A2(_02625_),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10509_ (.A1(_02767_),
    .A2(_02768_),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10510_ (.I(_02540_),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10511_ (.A1(_01552_),
    .A2(_02541_),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10512_ (.I(_02543_),
    .Z(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10513_ (.I(_02388_),
    .Z(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10514_ (.A1(_01679_),
    .A2(_02773_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10515_ (.A1(_01560_),
    .A2(_02772_),
    .B(_02774_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10516_ (.I(_02501_),
    .Z(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10517_ (.A1(_02770_),
    .A2(_02771_),
    .B(_02775_),
    .C(_02776_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10518_ (.I(_02777_),
    .Z(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10519_ (.I(_02778_),
    .Z(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10520_ (.A1(_02506_),
    .A2(_02779_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10521_ (.A1(_02769_),
    .A2(_02780_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10522_ (.A1(_02765_),
    .A2(_02781_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10523_ (.A1(_02743_),
    .A2(_02782_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10524_ (.A1(_02740_),
    .A2(_02783_),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _10525_ (.A1(_02735_),
    .A2(_02738_),
    .A3(_02784_),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10526_ (.I(_01100_),
    .Z(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10527_ (.A1(\channels.sample3[0] ),
    .A2(_02786_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10528_ (.A1(_02361_),
    .A2(_02785_),
    .B(_02787_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10529_ (.A1(_02738_),
    .A2(_02784_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10530_ (.A1(_02738_),
    .A2(_02784_),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10531_ (.A1(_02735_),
    .A2(_02788_),
    .B(_02789_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10532_ (.A1(_02743_),
    .A2(_02782_),
    .Z(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10533_ (.A1(_02740_),
    .A2(_02783_),
    .B(_02791_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10534_ (.A1(_02688_),
    .A2(_02626_),
    .A3(_02767_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10535_ (.A1(_02769_),
    .A2(_02780_),
    .B(_02793_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10536_ (.A1(_02746_),
    .A2(_02764_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10537_ (.A1(_02765_),
    .A2(_02781_),
    .B(_02795_),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10538_ (.A1(_02749_),
    .A2(_02756_),
    .Z(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10539_ (.A1(_02749_),
    .A2(_02756_),
    .Z(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10540_ (.A1(_02797_),
    .A2(_02763_),
    .B(_02798_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10541_ (.A1(_02750_),
    .A2(_02751_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10542_ (.A1(_02750_),
    .A2(_02751_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10543_ (.A1(_02800_),
    .A2(_02755_),
    .B(_02801_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10544_ (.A1(_02531_),
    .A2(_02636_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10545_ (.A1(_01167_),
    .A2(_02637_),
    .B(_02803_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10546_ (.A1(_02714_),
    .A2(_02804_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10547_ (.A1(_01698_),
    .A2(_02574_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10548_ (.A1(_02531_),
    .A2(_02575_),
    .B(_02806_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10549_ (.A1(_02752_),
    .A2(_02807_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10550_ (.A1(_02585_),
    .A2(_02592_),
    .Z(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10551_ (.A1(_02805_),
    .A2(_02808_),
    .A3(_02809_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10552_ (.A1(_02802_),
    .A2(_02810_),
    .Z(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10553_ (.A1(_02524_),
    .A2(_02624_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10554_ (.A1(_02546_),
    .A2(_02556_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10555_ (.A1(_02537_),
    .A2(_02502_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10556_ (.A1(_02813_),
    .A2(_02814_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10557_ (.A1(_02812_),
    .A2(_02815_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10558_ (.A1(_02811_),
    .A2(_02816_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10559_ (.A1(_02799_),
    .A2(_02817_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10560_ (.A1(_02757_),
    .A2(_02762_),
    .B(_02760_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10561_ (.A1(_02563_),
    .A2(_02778_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10562_ (.A1(_02819_),
    .A2(_02820_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10563_ (.A1(_01560_),
    .A2(_02569_),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10564_ (.A1(_01700_),
    .A2(_02773_),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10565_ (.A1(_01566_),
    .A2(_02772_),
    .B(_02823_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10566_ (.A1(_02770_),
    .A2(_02822_),
    .B(_02824_),
    .C(_02776_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10567_ (.I(_02825_),
    .Z(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10568_ (.A1(_02609_),
    .A2(_02826_),
    .ZN(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10569_ (.A1(_02821_),
    .A2(_02827_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10570_ (.A1(_02818_),
    .A2(_02828_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10571_ (.A1(_02796_),
    .A2(_02829_),
    .Z(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10572_ (.A1(_02794_),
    .A2(_02830_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10573_ (.A1(_02792_),
    .A2(_02831_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10574_ (.A1(_02790_),
    .A2(_02832_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10575_ (.A1(\channels.sample3[1] ),
    .A2(_02786_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10576_ (.A1(_02361_),
    .A2(_02833_),
    .B(_02834_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10577_ (.I(_02832_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10578_ (.A1(_02792_),
    .A2(_02831_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10579_ (.A1(_02790_),
    .A2(_02835_),
    .B(_02836_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10580_ (.A1(_02796_),
    .A2(_02829_),
    .Z(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10581_ (.A1(_02794_),
    .A2(_02830_),
    .B(_02838_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10582_ (.A1(_02689_),
    .A2(_02779_),
    .A3(_02819_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10583_ (.I(_02705_),
    .Z(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10584_ (.I(_02826_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10585_ (.A1(_02841_),
    .A2(_02821_),
    .A3(_02842_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10586_ (.A1(_02840_),
    .A2(_02843_),
    .Z(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10587_ (.A1(_02799_),
    .A2(_02817_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10588_ (.A1(_02818_),
    .A2(_02828_),
    .B(_02845_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10589_ (.A1(_02802_),
    .A2(_02810_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10590_ (.A1(_02811_),
    .A2(_02816_),
    .B(_02847_),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10591_ (.I(_02804_),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10592_ (.A1(_02752_),
    .A2(_02807_),
    .B1(_02849_),
    .B2(_02715_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10593_ (.A1(_02715_),
    .A2(_02752_),
    .A3(_02807_),
    .A4(_02849_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10594_ (.A1(_02850_),
    .A2(_02809_),
    .B(_02851_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10595_ (.A1(_02556_),
    .A2(_02603_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10596_ (.A1(_02510_),
    .A2(_02515_),
    .A3(_02639_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10597_ (.A1(_02577_),
    .A2(_02591_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10598_ (.A1(_02854_),
    .A2(_02855_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10599_ (.A1(_02853_),
    .A2(_02856_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10600_ (.A1(_02852_),
    .A2(_02857_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10601_ (.A1(_02852_),
    .A2(_02857_),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10602_ (.A1(_02858_),
    .A2(_02859_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10603_ (.A1(_02643_),
    .A2(_02777_),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10604_ (.A1(_02596_),
    .A2(_02502_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10605_ (.A1(_02538_),
    .A2(_02624_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10606_ (.A1(_02862_),
    .A2(_02863_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10607_ (.A1(_02861_),
    .A2(_02864_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10608_ (.A1(_02860_),
    .A2(_02865_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10609_ (.A1(_02813_),
    .A2(_02814_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10610_ (.A1(_02812_),
    .A2(_02815_),
    .B(_02867_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10611_ (.A1(_02564_),
    .A2(_02825_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10612_ (.A1(_02868_),
    .A2(_02869_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10613_ (.A1(_01566_),
    .A2(_02569_),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10614_ (.A1(_01716_),
    .A2(_02773_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10615_ (.A1(_02404_),
    .A2(_02772_),
    .B(_02872_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10616_ (.A1(_02770_),
    .A2(_02871_),
    .B(_02873_),
    .C(_02776_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10617_ (.I(_02874_),
    .Z(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10618_ (.A1(_02506_),
    .A2(_02875_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10619_ (.A1(_02870_),
    .A2(_02876_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10620_ (.A1(_02848_),
    .A2(_02866_),
    .A3(_02877_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10621_ (.A1(_02846_),
    .A2(_02878_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10622_ (.A1(_02844_),
    .A2(_02879_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10623_ (.A1(_02839_),
    .A2(_02880_),
    .Z(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10624_ (.A1(_02837_),
    .A2(_02881_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10625_ (.A1(\channels.sample3[2] ),
    .A2(_02786_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10626_ (.A1(_02361_),
    .A2(_02882_),
    .B(_02883_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10627_ (.I(_02360_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10628_ (.I(_02881_),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10629_ (.A1(_02839_),
    .A2(_02880_),
    .Z(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10630_ (.A1(_02837_),
    .A2(_02885_),
    .B(_02886_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10631_ (.A1(_02846_),
    .A2(_02878_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10632_ (.A1(_02844_),
    .A2(_02879_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10633_ (.A1(_02888_),
    .A2(_02889_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10634_ (.A1(_02689_),
    .A2(_02842_),
    .A3(_02868_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10635_ (.I(_02875_),
    .Z(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10636_ (.A1(_02841_),
    .A2(_02870_),
    .A3(_02892_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10637_ (.A1(_02891_),
    .A2(_02893_),
    .Z(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10638_ (.A1(_02848_),
    .A2(_02866_),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10639_ (.A1(_02848_),
    .A2(_02866_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10640_ (.A1(_02895_),
    .A2(_02877_),
    .B(_02896_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10641_ (.A1(_02860_),
    .A2(_02865_),
    .B(_02858_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10642_ (.A1(_02854_),
    .A2(_02855_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10643_ (.A1(_02853_),
    .A2(_02856_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10644_ (.A1(_02899_),
    .A2(_02900_),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10645_ (.A1(_02503_),
    .A2(_02603_),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10646_ (.A1(_02592_),
    .A2(_02639_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10647_ (.A1(_02555_),
    .A2(_02577_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10648_ (.A1(_02903_),
    .A2(_02904_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10649_ (.A1(_02902_),
    .A2(_02905_),
    .Z(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10650_ (.A1(_02902_),
    .A2(_02905_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10651_ (.A1(_02906_),
    .A2(_02907_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10652_ (.A1(_02901_),
    .A2(_02908_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10653_ (.A1(_02644_),
    .A2(_02825_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10654_ (.A1(_02659_),
    .A2(_02624_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10655_ (.A1(_02646_),
    .A2(_02777_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10656_ (.A1(_02911_),
    .A2(_02912_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10657_ (.A1(_02910_),
    .A2(_02913_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10658_ (.A1(_02909_),
    .A2(_02914_),
    .Z(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10659_ (.A1(_02898_),
    .A2(_02915_),
    .Z(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10660_ (.A1(_02862_),
    .A2(_02863_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10661_ (.A1(_02861_),
    .A2(_02864_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10662_ (.A1(_02917_),
    .A2(_02918_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10663_ (.A1(_02664_),
    .A2(_02874_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10664_ (.A1(_02919_),
    .A2(_02920_),
    .Z(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10665_ (.A1(_02404_),
    .A2(_02569_),
    .Z(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10666_ (.A1(_01726_),
    .A2(_02773_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10667_ (.A1(_01096_),
    .A2(_02772_),
    .B(_02923_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10668_ (.A1(_02770_),
    .A2(_02922_),
    .B(_02924_),
    .C(_02776_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10669_ (.A1(_02507_),
    .A2(_02925_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10670_ (.A1(_02921_),
    .A2(_02926_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10671_ (.A1(_02916_),
    .A2(_02927_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10672_ (.A1(_02897_),
    .A2(_02928_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10673_ (.A1(_02894_),
    .A2(_02929_),
    .Z(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10674_ (.A1(_02894_),
    .A2(_02929_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10675_ (.A1(_02930_),
    .A2(_02931_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10676_ (.A1(_02890_),
    .A2(_02932_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10677_ (.A1(_02887_),
    .A2(_02933_),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10678_ (.A1(\channels.sample3[3] ),
    .A2(_02786_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10679_ (.A1(_02884_),
    .A2(_02934_),
    .B(_02935_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10680_ (.I(_02933_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10681_ (.A1(_02890_),
    .A2(_02932_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10682_ (.A1(_02887_),
    .A2(_02936_),
    .B(_02937_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10683_ (.A1(_02897_),
    .A2(_02928_),
    .B(_02930_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10684_ (.A1(_02919_),
    .A2(_02920_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10685_ (.I(_02925_),
    .Z(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10686_ (.I(_02941_),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10687_ (.A1(_02841_),
    .A2(_02921_),
    .A3(_02942_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10688_ (.A1(_02940_),
    .A2(_02943_),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10689_ (.A1(_02898_),
    .A2(_02915_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10690_ (.A1(_02916_),
    .A2(_02927_),
    .B(_02945_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10691_ (.A1(_02911_),
    .A2(_02912_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10692_ (.A1(_02910_),
    .A2(_02913_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10693_ (.A1(_02947_),
    .A2(_02948_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10694_ (.A1(_02688_),
    .A2(_02925_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10695_ (.A1(_02949_),
    .A2(_02950_),
    .Z(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10696_ (.A1(_02901_),
    .A2(_02908_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10697_ (.A1(_02909_),
    .A2(_02914_),
    .B(_02952_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10698_ (.A1(_02903_),
    .A2(_02904_),
    .B(_02906_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10699_ (.A1(_02604_),
    .A2(_02625_),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10700_ (.A1(_02557_),
    .A2(_02640_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10701_ (.I(_02578_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10702_ (.A1(_02503_),
    .A2(_02957_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10703_ (.A1(_02956_),
    .A2(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10704_ (.A1(_02955_),
    .A2(_02959_),
    .Z(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10705_ (.A1(_02954_),
    .A2(_02960_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10706_ (.A1(_02712_),
    .A2(_02875_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10707_ (.I(_02659_),
    .Z(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10708_ (.A1(_02963_),
    .A2(_02779_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10709_ (.A1(_02678_),
    .A2(_02826_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10710_ (.A1(_02964_),
    .A2(_02965_),
    .Z(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10711_ (.A1(_02964_),
    .A2(_02965_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10712_ (.A1(_02966_),
    .A2(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10713_ (.A1(_02962_),
    .A2(_02968_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10714_ (.A1(_02961_),
    .A2(_02969_),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10715_ (.A1(_02951_),
    .A2(_02953_),
    .A3(_02970_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10716_ (.A1(_02946_),
    .A2(_02971_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10717_ (.A1(_02944_),
    .A2(_02972_),
    .Z(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10718_ (.A1(_02939_),
    .A2(_02973_),
    .Z(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10719_ (.A1(_02938_),
    .A2(_02974_),
    .Z(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10720_ (.I(_01099_),
    .Z(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10721_ (.I(_02976_),
    .Z(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10722_ (.A1(\channels.sample3[4] ),
    .A2(_02977_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10723_ (.A1(_02884_),
    .A2(_02975_),
    .B(_02978_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10724_ (.I(_02974_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10725_ (.A1(_02939_),
    .A2(_02973_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10726_ (.A1(_02938_),
    .A2(_02979_),
    .B(_02980_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10727_ (.A1(_02946_),
    .A2(_02971_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10728_ (.A1(_02944_),
    .A2(_02972_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10729_ (.A1(_02982_),
    .A2(_02983_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10730_ (.A1(_02949_),
    .A2(_02950_),
    .Z(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10731_ (.A1(_02953_),
    .A2(_02970_),
    .Z(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10732_ (.A1(_02953_),
    .A2(_02970_),
    .Z(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10733_ (.A1(_02951_),
    .A2(_02986_),
    .B(_02987_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10734_ (.A1(_02962_),
    .A2(_02968_),
    .B(_02966_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10735_ (.A1(_02954_),
    .A2(_02960_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10736_ (.A1(_02961_),
    .A2(_02969_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10737_ (.A1(_02990_),
    .A2(_02991_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10738_ (.A1(_02955_),
    .A2(_02959_),
    .Z(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10739_ (.A1(_02956_),
    .A2(_02958_),
    .B(_02993_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10740_ (.A1(_02604_),
    .A2(_02778_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10741_ (.I(_02640_),
    .Z(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10742_ (.A1(_02504_),
    .A2(_02996_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10743_ (.A1(_02957_),
    .A2(_02625_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10744_ (.A1(_02997_),
    .A2(_02998_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10745_ (.A1(_02995_),
    .A2(_02999_),
    .Z(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10746_ (.A1(_02994_),
    .A2(_03000_),
    .Z(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10747_ (.A1(_02712_),
    .A2(_02925_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10748_ (.A1(_02659_),
    .A2(_02825_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10749_ (.A1(_02678_),
    .A2(_02874_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10750_ (.A1(_03003_),
    .A2(_03004_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10751_ (.A1(_03002_),
    .A2(_03005_),
    .Z(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10752_ (.A1(_03001_),
    .A2(_03006_),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10753_ (.A1(_02992_),
    .A2(_03007_),
    .Z(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10754_ (.A1(_02989_),
    .A2(_03008_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10755_ (.A1(_02988_),
    .A2(_03009_),
    .Z(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10756_ (.A1(_02988_),
    .A2(_03009_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10757_ (.A1(_03010_),
    .A2(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10758_ (.A1(_02985_),
    .A2(_03012_),
    .Z(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10759_ (.A1(_02984_),
    .A2(_03013_),
    .Z(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10760_ (.A1(_02981_),
    .A2(_03014_),
    .Z(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10761_ (.A1(_01939_),
    .A2(_02977_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10762_ (.A1(_02884_),
    .A2(_03015_),
    .B(_03016_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10763_ (.A1(_02982_),
    .A2(_02983_),
    .B(_03013_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10764_ (.I(_03014_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10765_ (.A1(_02981_),
    .A2(_03018_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10766_ (.A1(_03017_),
    .A2(_03019_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10767_ (.A1(_02992_),
    .A2(_03007_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10768_ (.A1(_02989_),
    .A2(_03008_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10769_ (.A1(_03003_),
    .A2(_03004_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10770_ (.A1(_03002_),
    .A2(_03005_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10771_ (.A1(_02994_),
    .A2(_03000_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10772_ (.A1(_03001_),
    .A2(_03006_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10773_ (.A1(_03025_),
    .A2(_03026_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10774_ (.A1(_02995_),
    .A2(_02999_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10775_ (.A1(_02997_),
    .A2(_02998_),
    .B(_03028_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10776_ (.I(_02604_),
    .Z(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10777_ (.A1(_03030_),
    .A2(_02842_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10778_ (.A1(_02626_),
    .A2(_02996_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10779_ (.I(_02957_),
    .Z(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10780_ (.A1(_03033_),
    .A2(_02779_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10781_ (.A1(_03032_),
    .A2(_03034_),
    .Z(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10782_ (.A1(_03032_),
    .A2(_03034_),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10783_ (.A1(_03035_),
    .A2(_03036_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10784_ (.A1(_03031_),
    .A2(_03037_),
    .Z(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10785_ (.A1(_03029_),
    .A2(_03038_),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10786_ (.A1(_02963_),
    .A2(_02875_),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10787_ (.I(_02678_),
    .Z(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10788_ (.A1(_03041_),
    .A2(_02941_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10789_ (.A1(_03040_),
    .A2(_03042_),
    .Z(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10790_ (.A1(_03039_),
    .A2(_03043_),
    .Z(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10791_ (.A1(_03027_),
    .A2(_03044_),
    .Z(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10792_ (.A1(_03023_),
    .A2(_03024_),
    .B(_03045_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10793_ (.A1(_03023_),
    .A2(_03024_),
    .A3(_03045_),
    .Z(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10794_ (.A1(_03046_),
    .A2(_03047_),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10795_ (.A1(_03021_),
    .A2(_03022_),
    .B(_03048_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10796_ (.A1(_03021_),
    .A2(_03022_),
    .A3(_03048_),
    .Z(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10797_ (.A1(_03049_),
    .A2(_03050_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10798_ (.A1(_02985_),
    .A2(_03012_),
    .B(_03010_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10799_ (.A1(_03051_),
    .A2(_03052_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10800_ (.A1(_03020_),
    .A2(_03053_),
    .Z(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10801_ (.A1(\channels.sample3[6] ),
    .A2(_02977_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10802_ (.A1(_02884_),
    .A2(_03054_),
    .B(_03055_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10803_ (.I(_02360_),
    .Z(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10804_ (.A1(_03051_),
    .A2(_03052_),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10805_ (.A1(_03017_),
    .A2(_03019_),
    .B(_03053_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10806_ (.A1(_03057_),
    .A2(_03058_),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10807_ (.A1(_03040_),
    .A2(_03042_),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10808_ (.A1(_03029_),
    .A2(_03038_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10809_ (.A1(_03039_),
    .A2(_03043_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10810_ (.A1(_03061_),
    .A2(_03062_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10811_ (.A1(_02963_),
    .A2(_02941_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10812_ (.A1(_03031_),
    .A2(_03037_),
    .B(_03035_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10813_ (.A1(_03030_),
    .A2(_02874_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10814_ (.A1(_02996_),
    .A2(_02778_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10815_ (.A1(_02957_),
    .A2(_02826_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10816_ (.A1(_03067_),
    .A2(_03068_),
    .Z(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10817_ (.A1(_03067_),
    .A2(_03068_),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10818_ (.A1(_03069_),
    .A2(_03070_),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10819_ (.A1(_03066_),
    .A2(_03071_),
    .Z(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10820_ (.A1(_03065_),
    .A2(_03072_),
    .Z(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10821_ (.A1(_03064_),
    .A2(_03073_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10822_ (.A1(_03063_),
    .A2(_03074_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10823_ (.A1(_03060_),
    .A2(_03075_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10824_ (.A1(_03027_),
    .A2(_03044_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10825_ (.A1(_03077_),
    .A2(_03046_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10826_ (.A1(_03076_),
    .A2(_03078_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10827_ (.A1(_03049_),
    .A2(_03079_),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10828_ (.I(_03080_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10829_ (.A1(_03059_),
    .A2(_03081_),
    .Z(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10830_ (.A1(_01989_),
    .A2(_02977_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10831_ (.A1(_03056_),
    .A2(_03082_),
    .B(_03083_),
    .ZN(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10832_ (.I(_03079_),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10833_ (.A1(_03049_),
    .A2(_03084_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10834_ (.A1(_03057_),
    .A2(_03058_),
    .B(_03081_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10835_ (.A1(_03085_),
    .A2(_03086_),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10836_ (.A1(_03076_),
    .A2(_03078_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10837_ (.A1(_03030_),
    .A2(_02941_),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10838_ (.I(_02996_),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10839_ (.A1(_03090_),
    .A2(_02842_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10840_ (.A1(_03033_),
    .A2(_02892_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10841_ (.A1(_03089_),
    .A2(_03091_),
    .A3(_03092_),
    .Z(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10842_ (.A1(_03066_),
    .A2(_03071_),
    .B(_03069_),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10843_ (.I(_03094_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10844_ (.A1(_03093_),
    .A2(_03095_),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10845_ (.A1(_03065_),
    .A2(_03072_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10846_ (.I(_02963_),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10847_ (.A1(_03098_),
    .A2(_02942_),
    .A3(_03073_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10848_ (.A1(_03097_),
    .A2(_03099_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10849_ (.A1(_03096_),
    .A2(_03100_),
    .Z(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10850_ (.A1(_03063_),
    .A2(_03074_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10851_ (.A1(_03060_),
    .A2(_03075_),
    .B(_03102_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10852_ (.A1(_03101_),
    .A2(_03103_),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10853_ (.A1(_03088_),
    .A2(_03104_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10854_ (.A1(_03087_),
    .A2(_03105_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10855_ (.I(_02976_),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10856_ (.A1(\channels.sample3[8] ),
    .A2(_03107_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10857_ (.A1(_03056_),
    .A2(_03106_),
    .B(_03108_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10858_ (.A1(_03088_),
    .A2(_03104_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10859_ (.A1(_03087_),
    .A2(_03105_),
    .B(_03109_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10860_ (.A1(_03101_),
    .A2(_03103_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10861_ (.A1(_03091_),
    .A2(_03092_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10862_ (.A1(_03091_),
    .A2(_03092_),
    .Z(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10863_ (.A1(_03089_),
    .A2(_03112_),
    .B(_03113_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10864_ (.A1(_03090_),
    .A2(_02892_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10865_ (.A1(_03033_),
    .A2(_02942_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10866_ (.A1(_03115_),
    .A2(_03116_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10867_ (.A1(_03114_),
    .A2(_03117_),
    .Z(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10868_ (.A1(_03093_),
    .A2(_03095_),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10869_ (.A1(_03096_),
    .A2(_03100_),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10870_ (.A1(_03119_),
    .A2(_03120_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10871_ (.A1(_03118_),
    .A2(_03121_),
    .Z(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10872_ (.A1(_03111_),
    .A2(_03122_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10873_ (.A1(_03110_),
    .A2(_03123_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10874_ (.A1(_02040_),
    .A2(_03107_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10875_ (.A1(_03056_),
    .A2(_03124_),
    .B(_03125_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10876_ (.A1(_03110_),
    .A2(_03123_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10877_ (.A1(_03111_),
    .A2(_03122_),
    .B(_03126_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10878_ (.A1(_03120_),
    .A2(_03118_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10879_ (.A1(_03119_),
    .A2(_03118_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10880_ (.I(_03033_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10881_ (.A1(_03114_),
    .A2(_03117_),
    .Z(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10882_ (.A1(_03130_),
    .A2(_02892_),
    .B(_03131_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10883_ (.I(_03090_),
    .Z(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10884_ (.A1(_03133_),
    .A2(_02942_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10885_ (.I0(_03132_),
    .I1(_03131_),
    .S(_03134_),
    .Z(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10886_ (.A1(_03129_),
    .A2(_03135_),
    .Z(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10887_ (.A1(_03128_),
    .A2(_03136_),
    .Z(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10888_ (.A1(_03127_),
    .A2(_03137_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10889_ (.A1(\channels.sample3[10] ),
    .A2(_03107_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10890_ (.A1(_03056_),
    .A2(_03138_),
    .B(_03139_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10891_ (.I(_02360_),
    .Z(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10892_ (.A1(_03129_),
    .A2(_03132_),
    .B(_03134_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10893_ (.A1(_03128_),
    .A2(_03136_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10894_ (.A1(_03127_),
    .A2(_03137_),
    .B(_03141_),
    .C(_03142_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10895_ (.A1(_02068_),
    .A2(_03107_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10896_ (.A1(_03140_),
    .A2(_03143_),
    .B(_03144_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10897_ (.I(_01114_),
    .Z(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10898_ (.A1(\channels.sample2[0] ),
    .A2(_03145_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10899_ (.A1(_02368_),
    .A2(_02785_),
    .B(_03146_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10900_ (.A1(\channels.sample2[1] ),
    .A2(_03145_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10901_ (.A1(_02368_),
    .A2(_02833_),
    .B(_03147_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10902_ (.A1(\channels.sample2[2] ),
    .A2(_03145_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10903_ (.A1(_02368_),
    .A2(_02882_),
    .B(_03148_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10904_ (.I(_02367_),
    .Z(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10905_ (.A1(\channels.sample2[3] ),
    .A2(_03145_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10906_ (.A1(_03149_),
    .A2(_02934_),
    .B(_03150_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10907_ (.I(_01113_),
    .Z(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10908_ (.I(_03151_),
    .Z(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10909_ (.A1(\channels.sample2[4] ),
    .A2(_03152_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10910_ (.A1(_03149_),
    .A2(_02975_),
    .B(_03153_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10911_ (.A1(\channels.sample2[5] ),
    .A2(_03152_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10912_ (.A1(_03149_),
    .A2(_03015_),
    .B(_03154_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10913_ (.A1(\channels.sample2[6] ),
    .A2(_03152_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10914_ (.A1(_03149_),
    .A2(_03054_),
    .B(_03155_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10915_ (.I(_02367_),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10916_ (.A1(\channels.sample2[7] ),
    .A2(_03152_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10917_ (.A1(_03156_),
    .A2(_03082_),
    .B(_03157_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10918_ (.I(_03151_),
    .Z(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10919_ (.A1(\channels.sample2[8] ),
    .A2(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10920_ (.A1(_03156_),
    .A2(_03106_),
    .B(_03159_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10921_ (.A1(\channels.sample2[9] ),
    .A2(_03158_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10922_ (.A1(_03156_),
    .A2(_03124_),
    .B(_03160_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10923_ (.A1(\channels.sample2[10] ),
    .A2(_03158_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10924_ (.A1(_03156_),
    .A2(_03138_),
    .B(_03161_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10925_ (.I(_02367_),
    .Z(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10926_ (.A1(\channels.sample2[11] ),
    .A2(_03158_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10927_ (.A1(_03162_),
    .A2(_03143_),
    .B(_03163_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10928_ (.I(_01331_),
    .Z(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10929_ (.A1(\channels.sample1[0] ),
    .A2(_01570_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10930_ (.A1(_03164_),
    .A2(_02785_),
    .B(_03165_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10931_ (.I(_01470_),
    .Z(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10932_ (.A1(\channels.sample1[1] ),
    .A2(_03166_),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10933_ (.A1(_03164_),
    .A2(_02833_),
    .B(_03167_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10934_ (.A1(\channels.sample1[2] ),
    .A2(_03166_),
    .ZN(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10935_ (.A1(_03164_),
    .A2(_02882_),
    .B(_03168_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10936_ (.A1(\channels.sample1[3] ),
    .A2(_03166_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10937_ (.A1(_03164_),
    .A2(_02934_),
    .B(_03169_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10938_ (.I(_01330_),
    .Z(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10939_ (.A1(\channels.sample1[4] ),
    .A2(_03166_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10940_ (.A1(_03170_),
    .A2(_02975_),
    .B(_03171_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10941_ (.I(_01470_),
    .Z(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10942_ (.A1(\channels.sample1[5] ),
    .A2(_03172_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10943_ (.A1(_03170_),
    .A2(_03015_),
    .B(_03173_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10944_ (.A1(\channels.sample1[6] ),
    .A2(_03172_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10945_ (.A1(_03170_),
    .A2(_03054_),
    .B(_03174_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10946_ (.A1(\channels.sample1[7] ),
    .A2(_03172_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10947_ (.A1(_03170_),
    .A2(_03082_),
    .B(_03175_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10948_ (.I(_01330_),
    .Z(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10949_ (.A1(\channels.sample1[8] ),
    .A2(_03172_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10950_ (.A1(_03176_),
    .A2(_03106_),
    .B(_03177_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10951_ (.A1(\channels.sample1[9] ),
    .A2(_01271_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10952_ (.A1(_03176_),
    .A2(_03124_),
    .B(_03178_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10953_ (.A1(\channels.sample1[10] ),
    .A2(_01271_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10954_ (.A1(_03176_),
    .A2(_03138_),
    .B(_03179_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10955_ (.A1(\channels.sample1[11] ),
    .A2(_01271_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10956_ (.A1(_03176_),
    .A2(_03143_),
    .B(_03180_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10957_ (.I(\filters.sample_filtered[0] ),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10958_ (.I(\filters.filter_step[2] ),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _10959_ (.I(_03182_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _10960_ (.I(\filters.filter_step[1] ),
    .Z(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10961_ (.I(_03184_),
    .Z(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10962_ (.I(\filters.filter_step[0] ),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10963_ (.A1(_03183_),
    .A2(_03185_),
    .A3(_03186_),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10964_ (.I(_03187_),
    .Z(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10965_ (.I(_03188_),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10966_ (.I(_03189_),
    .Z(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10967_ (.I(_03190_),
    .Z(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10968_ (.I(_03182_),
    .Z(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10969_ (.I(_03192_),
    .Z(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _10970_ (.I(\filters.filter_step[1] ),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10971_ (.I(_03194_),
    .Z(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10972_ (.I(_03195_),
    .Z(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10973_ (.I(\filters.filter_step[0] ),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10974_ (.I(_03197_),
    .Z(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10975_ (.I(_03198_),
    .Z(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10976_ (.I(\filters.band[0] ),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _10977_ (.A1(_03193_),
    .A2(_03196_),
    .A3(_03199_),
    .B(_03200_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10978_ (.I(_03201_),
    .Z(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10979_ (.I(_03199_),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10980_ (.I(_03193_),
    .Z(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10981_ (.I(_03185_),
    .Z(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10982_ (.I(_03205_),
    .Z(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10983_ (.A1(_03204_),
    .A2(_03206_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10984_ (.A1(_03203_),
    .A2(_03207_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10985_ (.I(_03208_),
    .Z(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10986_ (.A1(\filters.low[0] ),
    .A2(_03191_),
    .B(_03202_),
    .C(_03209_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10987_ (.A1(_03203_),
    .A2(_03207_),
    .Z(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10988_ (.I(_03211_),
    .Z(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10989_ (.A1(\filters.high[0] ),
    .A2(_03212_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10990_ (.A1(_03181_),
    .A2(_03210_),
    .A3(_03213_),
    .Z(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10991_ (.A1(_03210_),
    .A2(_03213_),
    .B(_03181_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10992_ (.I(_03206_),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10993_ (.I(_03203_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10994_ (.I(_03217_),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10995_ (.I(_03191_),
    .Z(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10996_ (.I(_03219_),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10997_ (.I(_03220_),
    .Z(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10998_ (.I(_03221_),
    .Z(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10999_ (.I(_03222_),
    .Z(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11000_ (.I(_03223_),
    .Z(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11001_ (.I(_03224_),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11002_ (.I(_03225_),
    .Z(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11003_ (.I(_03226_),
    .Z(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11004_ (.I(_03227_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11005_ (.A1(\filters.lp ),
    .A2(_03228_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11006_ (.I(_03209_),
    .Z(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11007_ (.I(_03230_),
    .Z(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11008_ (.I(_03231_),
    .Z(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11009_ (.I(_03232_),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11010_ (.I(_03233_),
    .Z(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11011_ (.I(_03234_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11012_ (.I(_03235_),
    .Z(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11013_ (.I(_03236_),
    .Z(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11014_ (.I(_03237_),
    .Z(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11015_ (.A1(_03206_),
    .A2(_03217_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11016_ (.I(_03183_),
    .Z(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11017_ (.I(_03240_),
    .Z(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11018_ (.A1(\filters.hp ),
    .A2(_03238_),
    .B1(_03239_),
    .B2(\filters.bp ),
    .C(_03241_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11019_ (.A1(_01080_),
    .A2(_03229_),
    .A3(_03242_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11020_ (.A1(_03216_),
    .A2(_03218_),
    .B(_03243_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11021_ (.I(_03244_),
    .Z(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11022_ (.I(_03243_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11023_ (.I(_03246_),
    .Z(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11024_ (.A1(_03214_),
    .A2(_03215_),
    .A3(_03245_),
    .B1(_03247_),
    .B2(_03181_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11025_ (.I(\filters.filter_step[2] ),
    .Z(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11026_ (.I(_03248_),
    .Z(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11027_ (.I(_03195_),
    .Z(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11028_ (.I(\filters.filter_step[0] ),
    .Z(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11029_ (.I(_03251_),
    .Z(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11030_ (.I(\filters.band[1] ),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11031_ (.A1(_03249_),
    .A2(_03250_),
    .A3(_03252_),
    .B(_03253_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11032_ (.I(_03254_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11033_ (.I(_03255_),
    .Z(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11034_ (.I(_03256_),
    .Z(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11035_ (.I(_03257_),
    .Z(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11036_ (.A1(\filters.low[1] ),
    .A2(_03190_),
    .B(_03258_),
    .C(_03208_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11037_ (.A1(\filters.high[1] ),
    .A2(_03211_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11038_ (.A1(_03259_),
    .A2(_03260_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11039_ (.A1(\filters.sample_filtered[1] ),
    .A2(_03261_),
    .Z(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11040_ (.A1(_03215_),
    .A2(_03262_),
    .Z(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11041_ (.A1(_03215_),
    .A2(_03262_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11042_ (.I(\filters.sample_filtered[1] ),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11043_ (.A1(_03245_),
    .A2(_03263_),
    .A3(_03264_),
    .B1(_03247_),
    .B2(_03265_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11044_ (.I(\filters.sample_filtered[2] ),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11045_ (.I(_03246_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11046_ (.I(_03244_),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11047_ (.A1(_03259_),
    .A2(_03260_),
    .B(_03265_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11048_ (.I(\filters.low[2] ),
    .Z(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11049_ (.I(\filters.band[2] ),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11050_ (.A1(_03192_),
    .A2(_03195_),
    .A3(_03198_),
    .B(_03271_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11051_ (.I(_03272_),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11052_ (.I(_03273_),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11053_ (.I(_03274_),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11054_ (.A1(_03270_),
    .A2(_03191_),
    .B(_03275_),
    .C(_03208_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11055_ (.A1(\filters.high[2] ),
    .A2(_03211_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11056_ (.A1(_03276_),
    .A2(_03277_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11057_ (.A1(\filters.sample_filtered[2] ),
    .A2(_03278_),
    .Z(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11058_ (.A1(_03269_),
    .A2(_03263_),
    .B(_03279_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11059_ (.A1(_03269_),
    .A2(_03263_),
    .A3(_03279_),
    .Z(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11060_ (.A1(_03280_),
    .A2(_03281_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11061_ (.A1(_03266_),
    .A2(_03267_),
    .B1(_03268_),
    .B2(_03282_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11062_ (.I(\filters.sample_filtered[3] ),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11063_ (.I(\filters.low[3] ),
    .Z(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11064_ (.I(_03194_),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11065_ (.I(\filters.band[3] ),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11066_ (.A1(_03248_),
    .A2(_03285_),
    .A3(_03251_),
    .B(_03286_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11067_ (.I(_03287_),
    .Z(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11068_ (.I(net69),
    .Z(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11069_ (.I(_03289_),
    .Z(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11070_ (.A1(_03284_),
    .A2(_03191_),
    .B(_03290_),
    .C(_03208_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11071_ (.A1(\filters.high[3] ),
    .A2(_03212_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11072_ (.A1(_03291_),
    .A2(_03292_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11073_ (.A1(\filters.sample_filtered[3] ),
    .A2(_03293_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11074_ (.I(_03294_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11075_ (.A1(\filters.sample_filtered[2] ),
    .A2(_03278_),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11076_ (.A1(_03296_),
    .A2(_03280_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11077_ (.A1(_03295_),
    .A2(_03297_),
    .Z(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11078_ (.A1(_03283_),
    .A2(_03267_),
    .B1(_03268_),
    .B2(_03298_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11079_ (.I(\filters.sample_filtered[4] ),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11080_ (.I(\filters.high[4] ),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11081_ (.I(\filters.band[4] ),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11082_ (.A1(_03248_),
    .A2(_03195_),
    .A3(_03251_),
    .B(_03301_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11083_ (.I(_03302_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11084_ (.I(_03303_),
    .Z(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11085_ (.A1(\filters.low[4] ),
    .A2(_03219_),
    .B(_03304_),
    .C(_03209_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11086_ (.A1(_03300_),
    .A2(_03209_),
    .B(_03305_),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11087_ (.A1(\filters.sample_filtered[4] ),
    .A2(_03306_),
    .Z(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11088_ (.A1(_03296_),
    .A2(_03280_),
    .B(_03295_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11089_ (.A1(\filters.sample_filtered[3] ),
    .A2(_03293_),
    .B(_03308_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11090_ (.A1(_03307_),
    .A2(_03309_),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11091_ (.A1(_03299_),
    .A2(_03267_),
    .B1(_03268_),
    .B2(_03310_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11092_ (.I(\filters.sample_filtered[5] ),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11093_ (.I(\filters.low[5] ),
    .Z(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11094_ (.I(_03182_),
    .Z(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11095_ (.I(_03285_),
    .Z(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11096_ (.I(_03197_),
    .Z(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11097_ (.I(\filters.band[5] ),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11098_ (.A1(_03313_),
    .A2(_03314_),
    .A3(_03315_),
    .B(_03316_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11099_ (.I(_03317_),
    .Z(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11100_ (.I(_03318_),
    .Z(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11101_ (.A1(_03312_),
    .A2(_03219_),
    .B(_03319_),
    .C(_03230_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11102_ (.A1(\filters.high[5] ),
    .A2(_03212_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11103_ (.A1(_03320_),
    .A2(_03321_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11104_ (.A1(\filters.sample_filtered[5] ),
    .A2(_03322_),
    .Z(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11105_ (.I(_03307_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11106_ (.A1(\filters.sample_filtered[4] ),
    .A2(_03306_),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11107_ (.A1(_03324_),
    .A2(_03309_),
    .B(_03325_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11108_ (.A1(_03323_),
    .A2(_03326_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11109_ (.A1(_03311_),
    .A2(_03267_),
    .B1(_03268_),
    .B2(_03327_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11110_ (.I(\filters.sample_filtered[6] ),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11111_ (.I(_03246_),
    .Z(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11112_ (.I(_03244_),
    .Z(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11113_ (.I(\filters.low[6] ),
    .Z(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11114_ (.I(\filters.band[6] ),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11115_ (.A1(_03249_),
    .A2(_03250_),
    .A3(_03252_),
    .B(_03332_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11116_ (.I(_03333_),
    .Z(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11117_ (.I(_03334_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11118_ (.A1(_03331_),
    .A2(_03220_),
    .B(_03335_),
    .C(_03230_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11119_ (.I(_03212_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11120_ (.A1(\filters.high[6] ),
    .A2(_03337_),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11121_ (.A1(_03336_),
    .A2(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11122_ (.A1(\filters.sample_filtered[6] ),
    .A2(_03339_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11123_ (.A1(_03320_),
    .A2(_03321_),
    .B(_03311_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11124_ (.A1(_03323_),
    .A2(_03326_),
    .B(_03341_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11125_ (.A1(_03340_),
    .A2(_03342_),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11126_ (.A1(_03328_),
    .A2(_03329_),
    .B1(_03330_),
    .B2(_03343_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11127_ (.I(\filters.sample_filtered[7] ),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11128_ (.I(\filters.high[7] ),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11129_ (.I(_03230_),
    .Z(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11130_ (.I(\filters.low[7] ),
    .Z(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11131_ (.I(_03220_),
    .Z(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _11132_ (.I(\filters.band[7] ),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11133_ (.A1(_03193_),
    .A2(_03250_),
    .A3(_03199_),
    .B(_03349_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11134_ (.I(_03350_),
    .Z(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11135_ (.I(_03351_),
    .Z(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11136_ (.A1(_03347_),
    .A2(_03348_),
    .B(_03352_),
    .C(_03231_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11137_ (.A1(_03345_),
    .A2(_03346_),
    .B(_03353_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11138_ (.A1(\filters.sample_filtered[7] ),
    .A2(_03354_),
    .Z(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11139_ (.I(_03340_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11140_ (.A1(_03356_),
    .A2(_03342_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11141_ (.A1(\filters.sample_filtered[6] ),
    .A2(_03339_),
    .B(_03357_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11142_ (.A1(_03355_),
    .A2(_03358_),
    .Z(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11143_ (.A1(_03344_),
    .A2(_03329_),
    .B1(_03330_),
    .B2(_03359_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11144_ (.I(\filters.sample_filtered[8] ),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11145_ (.I(\filters.high[8] ),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11146_ (.I(\filters.low[8] ),
    .Z(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11147_ (.I(\filters.band[8] ),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11148_ (.A1(_03193_),
    .A2(_03250_),
    .A3(_03199_),
    .B(_03363_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11149_ (.I(_03364_),
    .Z(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11150_ (.I(_03365_),
    .Z(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11151_ (.A1(_03362_),
    .A2(_03222_),
    .B(_03366_),
    .C(_03346_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11152_ (.A1(_03361_),
    .A2(_03232_),
    .B(_03367_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11153_ (.A1(\filters.sample_filtered[8] ),
    .A2(_03368_),
    .Z(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11154_ (.I(_03355_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11155_ (.A1(_03370_),
    .A2(_03358_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11156_ (.A1(\filters.sample_filtered[7] ),
    .A2(_03354_),
    .B(_03371_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11157_ (.A1(_03369_),
    .A2(_03372_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11158_ (.A1(_03360_),
    .A2(_03329_),
    .B1(_03330_),
    .B2(_03373_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11159_ (.I(\filters.sample_filtered[9] ),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11160_ (.I(\filters.high[9] ),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11161_ (.I(\filters.low[9] ),
    .Z(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11162_ (.I(_03219_),
    .Z(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11163_ (.I(_03377_),
    .Z(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11164_ (.I(_03378_),
    .Z(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11165_ (.I(_03379_),
    .Z(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11166_ (.I(_03285_),
    .Z(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11167_ (.I(\filters.band[9] ),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11168_ (.A1(_03249_),
    .A2(_03381_),
    .A3(_03252_),
    .B(_03382_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11169_ (.I(_03383_),
    .Z(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11170_ (.I(_03384_),
    .Z(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11171_ (.A1(_03376_),
    .A2(_03380_),
    .B(_03385_),
    .C(_03232_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11172_ (.A1(_03375_),
    .A2(_03233_),
    .B(_03386_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11173_ (.A1(\filters.sample_filtered[9] ),
    .A2(_03387_),
    .Z(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11174_ (.I(_03369_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11175_ (.A1(_03389_),
    .A2(_03372_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11176_ (.A1(\filters.sample_filtered[8] ),
    .A2(_03368_),
    .B(_03390_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11177_ (.A1(_03388_),
    .A2(_03391_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11178_ (.A1(_03374_),
    .A2(_03329_),
    .B1(_03330_),
    .B2(_03392_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11179_ (.I(\filters.sample_filtered[10] ),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11180_ (.I(_03246_),
    .Z(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11181_ (.I(_03244_),
    .Z(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11182_ (.I(\filters.low[10] ),
    .Z(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11183_ (.I(_03223_),
    .Z(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11184_ (.I(\filters.band[10] ),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11185_ (.A1(_03249_),
    .A2(_03381_),
    .A3(_03252_),
    .B(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11186_ (.I(_03399_),
    .Z(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11187_ (.A1(_03396_),
    .A2(_03397_),
    .B(_03400_),
    .C(_03234_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11188_ (.I(_03337_),
    .Z(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11189_ (.I(_03402_),
    .Z(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11190_ (.A1(\filters.high[10] ),
    .A2(_03403_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11191_ (.A1(_03401_),
    .A2(_03404_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11192_ (.A1(\filters.sample_filtered[10] ),
    .A2(_03405_),
    .Z(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11193_ (.I(_03388_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11194_ (.A1(_03407_),
    .A2(_03391_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11195_ (.A1(\filters.sample_filtered[9] ),
    .A2(_03387_),
    .B(_03408_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11196_ (.A1(_03406_),
    .A2(_03409_),
    .Z(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11197_ (.A1(_03393_),
    .A2(_03394_),
    .B1(_03395_),
    .B2(_03410_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11198_ (.I(\filters.sample_filtered[11] ),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11199_ (.I(\filters.high[11] ),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11200_ (.I(\filters.low[11] ),
    .Z(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11201_ (.I(\filters.band[11] ),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _11202_ (.A1(_03313_),
    .A2(_03381_),
    .A3(_03315_),
    .B(_03414_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11203_ (.A1(_03413_),
    .A2(_03225_),
    .B(_03415_),
    .C(_03235_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11204_ (.A1(_03412_),
    .A2(_03235_),
    .B(_03416_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11205_ (.A1(\filters.sample_filtered[11] ),
    .A2(_03417_),
    .Z(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11206_ (.I(_03406_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11207_ (.A1(_03419_),
    .A2(_03409_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11208_ (.A1(\filters.sample_filtered[10] ),
    .A2(_03405_),
    .B(_03420_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11209_ (.A1(_03418_),
    .A2(_03421_),
    .Z(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11210_ (.A1(_03411_),
    .A2(_03394_),
    .B1(_03395_),
    .B2(_03422_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11211_ (.I(\filters.sample_filtered[12] ),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11212_ (.I(\filters.low[12] ),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11213_ (.I(\filters.band[12] ),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11214_ (.I(_03397_),
    .Z(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11215_ (.A1(_03425_),
    .A2(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11216_ (.A1(_03424_),
    .A2(_03226_),
    .B(_03427_),
    .C(_03236_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11217_ (.I(_03403_),
    .Z(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11218_ (.I(_03429_),
    .Z(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11219_ (.A1(\filters.high[12] ),
    .A2(_03430_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11220_ (.A1(_03428_),
    .A2(_03431_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11221_ (.A1(\filters.sample_filtered[12] ),
    .A2(_03432_),
    .Z(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11222_ (.I(_03418_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11223_ (.A1(_03434_),
    .A2(_03421_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11224_ (.A1(\filters.sample_filtered[11] ),
    .A2(_03417_),
    .B(_03435_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11225_ (.A1(_03433_),
    .A2(_03436_),
    .Z(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11226_ (.A1(_03423_),
    .A2(_03394_),
    .B1(_03395_),
    .B2(_03437_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11227_ (.A1(_03428_),
    .A2(_03431_),
    .B(_03423_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11228_ (.I(_03433_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11229_ (.A1(_03439_),
    .A2(_03436_),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11230_ (.I(\filters.low[13] ),
    .Z(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11231_ (.I(\filters.band[13] ),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11232_ (.A1(_03442_),
    .A2(_03226_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11233_ (.A1(_03441_),
    .A2(_03227_),
    .B(_03443_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11234_ (.A1(\filters.high[13] ),
    .A2(_03237_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11235_ (.A1(_03237_),
    .A2(_03444_),
    .B(_03445_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11236_ (.A1(\filters.sample_filtered[13] ),
    .A2(_03446_),
    .Z(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11237_ (.A1(_03438_),
    .A2(_03440_),
    .A3(_03447_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11238_ (.I(_03447_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11239_ (.A1(_03438_),
    .A2(_03440_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11240_ (.A1(_03449_),
    .A2(_03450_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11241_ (.I(\filters.sample_filtered[13] ),
    .Z(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11242_ (.I(_03452_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11243_ (.A1(_03245_),
    .A2(_03448_),
    .A3(_03451_),
    .B1(_03247_),
    .B2(_03453_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11244_ (.I(\filters.sample_filtered[14] ),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11245_ (.I(_03454_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11246_ (.A1(_03452_),
    .A2(_03446_),
    .B(_03451_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11247_ (.I(\filters.low[14] ),
    .Z(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _11248_ (.I(\filters.band[14] ),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11249_ (.A1(_03458_),
    .A2(_03227_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11250_ (.A1(_03457_),
    .A2(_03228_),
    .B(_03459_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11251_ (.A1(\filters.high[14] ),
    .A2(_03237_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11252_ (.A1(_03238_),
    .A2(_03460_),
    .B(_03461_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11253_ (.A1(_03454_),
    .A2(_03462_),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11254_ (.A1(_03456_),
    .A2(_03463_),
    .Z(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11255_ (.A1(_03455_),
    .A2(_03394_),
    .B1(_03395_),
    .B2(_03464_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11256_ (.I(_03463_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11257_ (.A1(_03456_),
    .A2(_03465_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11258_ (.A1(_03454_),
    .A2(_03462_),
    .B(_03466_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11259_ (.I(\filters.sample_filtered[15] ),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11260_ (.I(\filters.high[15] ),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11261_ (.I(\filters.low[15] ),
    .Z(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11262_ (.A1(_03470_),
    .A2(_03228_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11263_ (.A1(_03204_),
    .A2(_03196_),
    .A3(_03203_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11264_ (.I(_03472_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11265_ (.I(_03473_),
    .Z(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11266_ (.I(_03474_),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11267_ (.I(_03475_),
    .Z(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11268_ (.I(_03476_),
    .Z(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11269_ (.I(_03477_),
    .Z(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11270_ (.I(_03478_),
    .Z(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11271_ (.A1(\filters.band[15] ),
    .A2(_03479_),
    .B(_03238_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _11272_ (.A1(_03469_),
    .A2(_03238_),
    .B1(_03471_),
    .B2(_03480_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11273_ (.A1(_03468_),
    .A2(_03481_),
    .Z(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11274_ (.A1(_03467_),
    .A2(_03482_),
    .Z(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11275_ (.A1(_03467_),
    .A2(_03482_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11276_ (.A1(_03245_),
    .A2(_03483_),
    .A3(_03484_),
    .B1(_03247_),
    .B2(_03468_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11277_ (.A1(_02100_),
    .A2(_01860_),
    .Z(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11278_ (.I(_03485_),
    .Z(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11279_ (.A1(\filters.cutoff_lut[6] ),
    .A2(_03486_),
    .B(_02345_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11280_ (.A1(_02309_),
    .A2(_03486_),
    .B(_03487_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11281_ (.I(_02337_),
    .Z(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11282_ (.A1(\filters.cutoff_lut[7] ),
    .A2(_03485_),
    .B(_03488_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11283_ (.A1(_02315_),
    .A2(_03486_),
    .B(_03489_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11284_ (.A1(\filters.cutoff_lut[8] ),
    .A2(_03485_),
    .B(_03488_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11285_ (.A1(_02318_),
    .A2(_03486_),
    .B(_03490_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11286_ (.I(\tt_um_rejunity_sn76489.control_tone_freq[0][0] ),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11287_ (.I(_01815_),
    .Z(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11288_ (.I(net12),
    .Z(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11289_ (.I(net11),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11290_ (.I(_03494_),
    .Z(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11291_ (.I(net14),
    .Z(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11292_ (.I(_01104_),
    .Z(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11293_ (.A1(_01829_),
    .A2(_01837_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _11294_ (.A1(_01835_),
    .A2(_01016_),
    .A3(_03498_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11295_ (.A1(_03497_),
    .A2(_03499_),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11296_ (.A1(_03496_),
    .A2(_03500_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11297_ (.I(_03501_),
    .Z(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11298_ (.A1(_03492_),
    .A2(_03493_),
    .A3(_03495_),
    .A4(_03502_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11299_ (.I(_03503_),
    .Z(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11300_ (.I(net7),
    .Z(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11301_ (.I(_03503_),
    .Z(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11302_ (.A1(_03505_),
    .A2(_03506_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11303_ (.I(_01760_),
    .Z(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11304_ (.I(_03508_),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11305_ (.I(_03509_),
    .Z(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11306_ (.A1(_03491_),
    .A2(_03504_),
    .B(_03507_),
    .C(_03510_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11307_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][1] ),
    .A2(_03506_),
    .B(_03488_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11308_ (.A1(_02315_),
    .A2(_03504_),
    .B(_03511_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11309_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][2] ),
    .A2(_03506_),
    .B(_03488_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11310_ (.A1(_02318_),
    .A2(_03504_),
    .B(_03512_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11311_ (.I(_02337_),
    .Z(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11312_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][3] ),
    .A2(_03506_),
    .B(_03513_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11313_ (.A1(_02321_),
    .A2(_03504_),
    .B(_03514_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11314_ (.I(\tt_um_rejunity_sn76489.control_tone_freq[2][0] ),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11315_ (.A1(_01816_),
    .A2(_03493_),
    .A3(_03495_),
    .A4(_03501_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11316_ (.I(_03516_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11317_ (.I(_03516_),
    .Z(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11318_ (.A1(_03505_),
    .A2(_03518_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11319_ (.A1(_03515_),
    .A2(_03517_),
    .B(_03519_),
    .C(_03510_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11320_ (.I(_02188_),
    .Z(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11321_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ),
    .A2(_03518_),
    .B(_03513_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11322_ (.A1(_03520_),
    .A2(_03517_),
    .B(_03521_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11323_ (.I(_02193_),
    .Z(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11324_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][2] ),
    .A2(_03518_),
    .B(_03513_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11325_ (.A1(_03522_),
    .A2(_03517_),
    .B(_03523_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11326_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][3] ),
    .A2(_03518_),
    .B(_03513_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11327_ (.A1(_02321_),
    .A2(_03517_),
    .B(_03524_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11328_ (.A1(_01810_),
    .A2(_03494_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11329_ (.A1(_01815_),
    .A2(_03501_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11330_ (.A1(_03525_),
    .A2(_03526_),
    .Z(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11331_ (.I(_03527_),
    .Z(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11332_ (.I(_03527_),
    .Z(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11333_ (.A1(_01750_),
    .A2(_03529_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11334_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][0] ),
    .A2(_03528_),
    .B(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11335_ (.A1(_03510_),
    .A2(_03531_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11336_ (.I(_02264_),
    .Z(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11337_ (.I(_03532_),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11338_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ),
    .A2(_03529_),
    .B(_03533_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11339_ (.A1(_03520_),
    .A2(_03528_),
    .B(_03534_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11340_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][2] ),
    .A2(_03529_),
    .B(_03533_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11341_ (.A1(_03522_),
    .A2(_03528_),
    .B(_03535_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11342_ (.I(_02320_),
    .Z(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11343_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][3] ),
    .A2(_03529_),
    .B(_03533_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11344_ (.A1(_03536_),
    .A2(_03528_),
    .B(_03537_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11345_ (.I0(\channels.adsr_state[0][0] ),
    .I1(\channels.adsr_state[1][0] ),
    .I2(\channels.adsr_state[2][0] ),
    .I3(\channels.adsr_state[3][0] ),
    .S0(_01156_),
    .S1(_01170_),
    .Z(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11346_ (.I(_03538_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11347_ (.I0(\channels.adsr_state[0][1] ),
    .I1(\channels.adsr_state[1][1] ),
    .I2(\channels.adsr_state[2][1] ),
    .I3(\channels.adsr_state[3][1] ),
    .S0(_01157_),
    .S1(_01171_),
    .Z(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11348_ (.A1(_03539_),
    .A2(_03540_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11349_ (.I(_03541_),
    .Z(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11350_ (.I(_03542_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11351_ (.I(_02807_),
    .Z(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11352_ (.I(_02712_),
    .Z(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11353_ (.A1(_02709_),
    .A2(_02713_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11354_ (.A1(_03041_),
    .A2(_03545_),
    .A3(_03546_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11355_ (.I(_03098_),
    .Z(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11356_ (.I(_03030_),
    .Z(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11357_ (.A1(_03548_),
    .A2(_03549_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11358_ (.A1(_03547_),
    .A2(_03550_),
    .Z(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11359_ (.A1(_03544_),
    .A2(_03551_),
    .Z(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11360_ (.A1(_02849_),
    .A2(_03552_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11361_ (.A1(_01595_),
    .A2(_03543_),
    .A3(_03553_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11362_ (.A1(_03543_),
    .A2(_03553_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11363_ (.A1(\channels.ctrl_reg2[0] ),
    .A2(_01292_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11364_ (.A1(\channels.ctrl_reg3[0] ),
    .A2(_01591_),
    .B1(_01305_),
    .B2(\channels.ctrl_reg1[0] ),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11365_ (.A1(_03556_),
    .A2(_03557_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11366_ (.A1(_03538_),
    .A2(_03540_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _11367_ (.A1(_03555_),
    .A2(_03558_),
    .A3(_03559_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11368_ (.I(_01052_),
    .Z(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11369_ (.A1(_01264_),
    .A2(_03560_),
    .B(_03561_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11370_ (.I0(_03554_),
    .I1(\channels.adsr_state[0][0] ),
    .S(_03562_),
    .Z(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11371_ (.I(_03563_),
    .Z(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11372_ (.A1(_01595_),
    .A2(_03538_),
    .A3(_03540_),
    .A4(_03558_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11373_ (.I0(_03564_),
    .I1(\channels.adsr_state[0][1] ),
    .S(_03562_),
    .Z(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11374_ (.I(_03565_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11375_ (.I(_01099_),
    .Z(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11376_ (.I(_03566_),
    .Z(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11377_ (.I(_01095_),
    .Z(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11378_ (.A1(_01321_),
    .A2(_03567_),
    .B1(_01326_),
    .B2(_03568_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11379_ (.I(_02976_),
    .Z(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11380_ (.A1(\channels.accum[2][1] ),
    .A2(_03569_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11381_ (.A1(_03140_),
    .A2(_01343_),
    .B(_03570_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11382_ (.I(\channels.accum[2][2] ),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11383_ (.A1(_03571_),
    .A2(_03567_),
    .B1(_01358_),
    .B2(_03568_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11384_ (.A1(\channels.accum[2][3] ),
    .A2(_03569_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11385_ (.A1(_03140_),
    .A2(_01369_),
    .B(_03572_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11386_ (.I(\channels.accum[2][4] ),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11387_ (.A1(_03573_),
    .A2(_03567_),
    .B1(_01382_),
    .B2(_03568_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11388_ (.A1(\channels.accum[2][5] ),
    .A2(_03569_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11389_ (.A1(_03140_),
    .A2(_01391_),
    .B(_03574_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11390_ (.I(\channels.accum[2][6] ),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11391_ (.A1(_03575_),
    .A2(_03567_),
    .B1(_01405_),
    .B2(_03568_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11392_ (.I(_02359_),
    .Z(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11393_ (.A1(\channels.accum[2][7] ),
    .A2(_03569_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11394_ (.A1(_03576_),
    .A2(_01416_),
    .B(_03577_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11395_ (.I(\channels.accum[2][8] ),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11396_ (.I(_01100_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11397_ (.I(_01250_),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11398_ (.A1(_03578_),
    .A2(_03579_),
    .B1(_01430_),
    .B2(_03580_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11399_ (.I(_02976_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11400_ (.A1(\channels.accum[2][9] ),
    .A2(_03581_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11401_ (.A1(_03576_),
    .A2(_01443_),
    .B(_03582_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11402_ (.I(\channels.accum[2][10] ),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11403_ (.A1(_03583_),
    .A2(_03579_),
    .B1(_01458_),
    .B2(_03580_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11404_ (.A1(\channels.accum[2][11] ),
    .A2(_03581_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11405_ (.A1(_03576_),
    .A2(_01469_),
    .B(_03584_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11406_ (.I(\channels.accum[2][12] ),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11407_ (.A1(_03585_),
    .A2(_03579_),
    .B1(_01485_),
    .B2(_03580_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11408_ (.A1(\channels.accum[2][13] ),
    .A2(_03581_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11409_ (.A1(_03576_),
    .A2(_01497_),
    .B(_03586_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11410_ (.I(\channels.accum[2][14] ),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11411_ (.A1(_03587_),
    .A2(_03579_),
    .B1(_01513_),
    .B2(_03580_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11412_ (.I(_02359_),
    .Z(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11413_ (.A1(\channels.accum[2][15] ),
    .A2(_03581_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11414_ (.A1(_03588_),
    .A2(_01525_),
    .B(_03589_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11415_ (.I(\channels.accum[2][16] ),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11416_ (.I(_01100_),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11417_ (.I(_01250_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11418_ (.A1(_03590_),
    .A2(_03591_),
    .B1(_01534_),
    .B2(_03592_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11419_ (.A1(\channels.accum[2][17] ),
    .A2(_01255_),
    .B1(_01540_),
    .B2(_01095_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11420_ (.I(_03593_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11421_ (.I(\channels.accum[2][18] ),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11422_ (.A1(_03594_),
    .A2(_03591_),
    .B1(_01549_),
    .B2(_03592_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11423_ (.A1(\channels.accum[2][19] ),
    .A2(_03566_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11424_ (.A1(_03588_),
    .A2(_01555_),
    .B(_03595_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11425_ (.I(\channels.accum[2][20] ),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11426_ (.A1(_03596_),
    .A2(_03591_),
    .B1(_01562_),
    .B2(_03592_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11427_ (.A1(\channels.accum[2][21] ),
    .A2(_03566_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11428_ (.A1(_03588_),
    .A2(_01569_),
    .B(_03597_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11429_ (.A1(_01574_),
    .A2(_03591_),
    .B1(_01578_),
    .B2(_03592_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11430_ (.A1(\channels.accum[2][23] ),
    .A2(_03566_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11431_ (.A1(_03588_),
    .A2(_01581_),
    .B(_03598_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11432_ (.I(\channels.accum[1][0] ),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11433_ (.I(_01113_),
    .Z(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11434_ (.I(_03600_),
    .Z(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11435_ (.I(_01112_),
    .Z(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11436_ (.A1(_03599_),
    .A2(_03601_),
    .B1(_01326_),
    .B2(_03602_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11437_ (.I(_03151_),
    .Z(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11438_ (.A1(\channels.accum[1][1] ),
    .A2(_03603_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11439_ (.A1(_03162_),
    .A2(_01343_),
    .B(_03604_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11440_ (.I(\channels.accum[1][2] ),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11441_ (.A1(_03605_),
    .A2(_03601_),
    .B1(_01358_),
    .B2(_03602_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11442_ (.A1(\channels.accum[1][3] ),
    .A2(_03603_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11443_ (.A1(_03162_),
    .A2(_01369_),
    .B(_03606_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11444_ (.I(\channels.accum[1][4] ),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11445_ (.A1(_03607_),
    .A2(_03601_),
    .B1(_01382_),
    .B2(_03602_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11446_ (.A1(\channels.accum[1][5] ),
    .A2(_03603_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11447_ (.A1(_03162_),
    .A2(_01391_),
    .B(_03608_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11448_ (.I(\channels.accum[1][6] ),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11449_ (.A1(_03609_),
    .A2(_03601_),
    .B1(_01405_),
    .B2(_03602_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11450_ (.I(_02366_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11451_ (.A1(\channels.accum[1][7] ),
    .A2(_03603_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11452_ (.A1(_03610_),
    .A2(_01416_),
    .B(_03611_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11453_ (.I(\channels.accum[1][8] ),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11454_ (.I(_01114_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11455_ (.I(_01229_),
    .Z(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11456_ (.A1(_03612_),
    .A2(_03613_),
    .B1(_01430_),
    .B2(_03614_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11457_ (.I(_03151_),
    .Z(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11458_ (.A1(\channels.accum[1][9] ),
    .A2(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11459_ (.A1(_03610_),
    .A2(_01443_),
    .B(_03616_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11460_ (.I(\channels.accum[1][10] ),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11461_ (.A1(_03617_),
    .A2(_03613_),
    .B1(_01458_),
    .B2(_03614_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11462_ (.A1(\channels.accum[1][11] ),
    .A2(_03615_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11463_ (.A1(_03610_),
    .A2(_01469_),
    .B(_03618_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11464_ (.I(\channels.accum[1][12] ),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11465_ (.A1(_03619_),
    .A2(_03613_),
    .B1(_01485_),
    .B2(_03614_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11466_ (.A1(\channels.accum[1][13] ),
    .A2(_03615_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11467_ (.A1(_03610_),
    .A2(_01497_),
    .B(_03620_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11468_ (.I(\channels.accum[1][14] ),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11469_ (.A1(_03621_),
    .A2(_03613_),
    .B1(_01513_),
    .B2(_03614_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11470_ (.I(_02366_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11471_ (.A1(\channels.accum[1][15] ),
    .A2(_03615_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11472_ (.A1(_03622_),
    .A2(_01525_),
    .B(_03623_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11473_ (.I(\channels.accum[1][16] ),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11474_ (.I(_01114_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11475_ (.I(_01229_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11476_ (.A1(_03624_),
    .A2(_03625_),
    .B1(_01534_),
    .B2(_03626_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11477_ (.A1(\channels.accum[1][17] ),
    .A2(_01240_),
    .B1(_01540_),
    .B2(_01112_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11478_ (.I(_03627_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11479_ (.I(\channels.accum[1][18] ),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11480_ (.A1(_03628_),
    .A2(_03625_),
    .B1(_01549_),
    .B2(_03626_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11481_ (.A1(\channels.accum[1][19] ),
    .A2(_03600_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11482_ (.A1(_03622_),
    .A2(_01555_),
    .B(_03629_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11483_ (.I(\channels.accum[1][20] ),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11484_ (.A1(_03630_),
    .A2(_03625_),
    .B1(_01562_),
    .B2(_03626_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11485_ (.A1(\channels.accum[1][21] ),
    .A2(_03600_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11486_ (.A1(_03622_),
    .A2(_01569_),
    .B(_03631_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11487_ (.A1(_01573_),
    .A2(_03625_),
    .B1(_01578_),
    .B2(_03626_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11488_ (.A1(\channels.accum[1][23] ),
    .A2(_03600_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11489_ (.A1(_03622_),
    .A2(_01581_),
    .B(_03632_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11490_ (.A1(_01037_),
    .A2(_01070_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11491_ (.I(_03633_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11492_ (.I(_00389_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11493_ (.A1(_02310_),
    .A2(_01966_),
    .Z(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11494_ (.I(_03634_),
    .Z(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11495_ (.I(_03635_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11496_ (.I(_03634_),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11497_ (.A1(\channels.freq1[0] ),
    .A2(_03637_),
    .B(_03533_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11498_ (.A1(_02309_),
    .A2(_03636_),
    .B(_03638_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11499_ (.I(_03532_),
    .Z(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11500_ (.A1(\channels.freq1[1] ),
    .A2(_03637_),
    .B(_03639_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11501_ (.A1(_03520_),
    .A2(_03636_),
    .B(_03640_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11502_ (.A1(\channels.freq1[2] ),
    .A2(_03637_),
    .B(_03639_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11503_ (.A1(_03522_),
    .A2(_03636_),
    .B(_03641_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11504_ (.A1(\channels.freq1[3] ),
    .A2(_03637_),
    .B(_03639_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11505_ (.A1(_03536_),
    .A2(_03636_),
    .B(_03642_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11506_ (.I(_02352_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11507_ (.A1(_03643_),
    .A2(_02023_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11508_ (.A1(\channels.freq1[4] ),
    .A2(_03644_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11509_ (.I(_03495_),
    .Z(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11510_ (.I(_03646_),
    .Z(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11511_ (.I(_03634_),
    .Z(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11512_ (.A1(_03647_),
    .A2(_03648_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11513_ (.I(_01098_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11514_ (.I(_03650_),
    .Z(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11515_ (.I(_03651_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11516_ (.A1(_03645_),
    .A2(_03649_),
    .B(_03652_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11517_ (.A1(\channels.freq1[5] ),
    .A2(_03635_),
    .B(_03639_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11518_ (.A1(_02326_),
    .A2(_03648_),
    .B(_03653_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11519_ (.I(_03532_),
    .Z(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11520_ (.A1(\channels.freq1[6] ),
    .A2(_03635_),
    .B(_03654_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11521_ (.A1(_02329_),
    .A2(_03648_),
    .B(_03655_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11522_ (.A1(\channels.freq1[7] ),
    .A2(_03635_),
    .B(_03654_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11523_ (.A1(_02331_),
    .A2(_03648_),
    .B(_03656_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11524_ (.I(_01750_),
    .Z(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11525_ (.I(_01789_),
    .Z(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11526_ (.A1(_03658_),
    .A2(_01894_),
    .Z(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11527_ (.I(_03659_),
    .Z(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11528_ (.I(_03660_),
    .Z(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11529_ (.I(_03660_),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11530_ (.A1(\channels.pw1[0] ),
    .A2(_03662_),
    .B(_03654_),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11531_ (.A1(_03657_),
    .A2(_03661_),
    .B(_03663_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11532_ (.I(_03659_),
    .Z(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11533_ (.A1(\channels.pw1[1] ),
    .A2(_03664_),
    .B(_03654_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11534_ (.A1(_03520_),
    .A2(_03661_),
    .B(_03665_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11535_ (.I(_03532_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11536_ (.A1(\channels.pw1[2] ),
    .A2(_03664_),
    .B(_03666_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11537_ (.A1(_03522_),
    .A2(_03661_),
    .B(_03667_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11538_ (.A1(\channels.pw1[3] ),
    .A2(_03664_),
    .B(_03666_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11539_ (.A1(_03536_),
    .A2(_03661_),
    .B(_03668_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11540_ (.A1(_02352_),
    .A2(_02015_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11541_ (.A1(_03646_),
    .A2(_03669_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11542_ (.I(_01827_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11543_ (.A1(_02441_),
    .A2(_03669_),
    .B(_03670_),
    .C(_03671_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11544_ (.A1(\channels.pw1[5] ),
    .A2(_03664_),
    .B(_03666_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11545_ (.A1(_02326_),
    .A2(_03662_),
    .B(_03672_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11546_ (.A1(\channels.pw1[6] ),
    .A2(_03660_),
    .B(_03666_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11547_ (.A1(_02329_),
    .A2(_03662_),
    .B(_03673_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11548_ (.I(_01071_),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11549_ (.I(_03674_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11550_ (.I(_03675_),
    .Z(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11551_ (.A1(\channels.pw1[7] ),
    .A2(_03660_),
    .B(_03676_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11552_ (.A1(_02331_),
    .A2(_03662_),
    .B(_03677_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11553_ (.A1(_02310_),
    .A2(_01890_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11554_ (.I(_03678_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11555_ (.I(_03679_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11556_ (.I(_03678_),
    .Z(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11557_ (.A1(\channels.freq2[0] ),
    .A2(_03681_),
    .B(_03676_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11558_ (.A1(_03657_),
    .A2(_03680_),
    .B(_03682_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11559_ (.I(_01765_),
    .Z(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11560_ (.A1(\channels.freq2[1] ),
    .A2(_03681_),
    .B(_03676_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11561_ (.A1(_03683_),
    .A2(_03680_),
    .B(_03684_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11562_ (.I(_01775_),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11563_ (.A1(\channels.freq2[2] ),
    .A2(_03681_),
    .B(_03676_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11564_ (.A1(_03685_),
    .A2(_03680_),
    .B(_03686_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11565_ (.I(_03675_),
    .Z(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11566_ (.A1(\channels.freq2[3] ),
    .A2(_03681_),
    .B(_03687_),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11567_ (.A1(_03536_),
    .A2(_03680_),
    .B(_03688_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11568_ (.A1(_03643_),
    .A2(_02013_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11569_ (.A1(\channels.freq2[4] ),
    .A2(_03689_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11570_ (.I(_03678_),
    .Z(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11571_ (.A1(_03647_),
    .A2(_03691_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11572_ (.A1(_03690_),
    .A2(_03692_),
    .B(_03652_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11573_ (.I(_02160_),
    .Z(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11574_ (.A1(\channels.freq2[5] ),
    .A2(_03679_),
    .B(_03687_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11575_ (.A1(_03693_),
    .A2(_03691_),
    .B(_03694_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11576_ (.I(_01816_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11577_ (.A1(\channels.freq2[6] ),
    .A2(_03679_),
    .B(_03687_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11578_ (.A1(_03695_),
    .A2(_03691_),
    .B(_03696_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11579_ (.I(_01821_),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11580_ (.A1(\channels.freq2[7] ),
    .A2(_03679_),
    .B(_03687_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11581_ (.A1(_03697_),
    .A2(_03691_),
    .B(_03698_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11582_ (.A1(_03658_),
    .A2(_01880_),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11583_ (.I(_03699_),
    .Z(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11584_ (.I(_03700_),
    .Z(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11585_ (.I(_03699_),
    .Z(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11586_ (.I(_03675_),
    .Z(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11587_ (.A1(\channels.freq3[0] ),
    .A2(_03702_),
    .B(_03703_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11588_ (.A1(_03657_),
    .A2(_03701_),
    .B(_03704_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11589_ (.A1(\channels.freq3[1] ),
    .A2(_03702_),
    .B(_03703_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11590_ (.A1(_03683_),
    .A2(_03701_),
    .B(_03705_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11591_ (.A1(\channels.freq3[2] ),
    .A2(_03702_),
    .B(_03703_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11592_ (.A1(_03685_),
    .A2(_03701_),
    .B(_03706_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11593_ (.I(_02320_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11594_ (.A1(\channels.freq3[3] ),
    .A2(_03702_),
    .B(_03703_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11595_ (.A1(_03707_),
    .A2(_03701_),
    .B(_03708_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11596_ (.A1(_03643_),
    .A2(_01949_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11597_ (.A1(\channels.freq3[4] ),
    .A2(_03709_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11598_ (.I(_03699_),
    .Z(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11599_ (.A1(_03647_),
    .A2(_03711_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11600_ (.A1(_03710_),
    .A2(_03712_),
    .B(_03652_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11601_ (.I(_03675_),
    .Z(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11602_ (.A1(\channels.freq3[5] ),
    .A2(_03700_),
    .B(_03713_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11603_ (.A1(_03693_),
    .A2(_03711_),
    .B(_03714_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11604_ (.A1(\channels.freq3[6] ),
    .A2(_03700_),
    .B(_03713_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11605_ (.A1(_03695_),
    .A2(_03711_),
    .B(_03715_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11606_ (.A1(\channels.freq3[7] ),
    .A2(_03700_),
    .B(_03713_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11607_ (.A1(_03697_),
    .A2(_03711_),
    .B(_03716_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11608_ (.A1(_03658_),
    .A2(_01907_),
    .Z(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11609_ (.I(_03717_),
    .Z(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11610_ (.I(_03718_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11611_ (.I(_03717_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11612_ (.A1(\channels.pw3[0] ),
    .A2(_03720_),
    .B(_03713_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11613_ (.A1(_03657_),
    .A2(_03719_),
    .B(_03721_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11614_ (.I(_03674_),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11615_ (.I(_03722_),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11616_ (.A1(\channels.pw3[1] ),
    .A2(_03720_),
    .B(_03723_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11617_ (.A1(_03683_),
    .A2(_03719_),
    .B(_03724_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11618_ (.A1(\channels.pw3[2] ),
    .A2(_03720_),
    .B(_03723_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11619_ (.A1(_03685_),
    .A2(_03719_),
    .B(_03725_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11620_ (.A1(\channels.pw3[3] ),
    .A2(_03720_),
    .B(_03723_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11621_ (.A1(_03707_),
    .A2(_03719_),
    .B(_03726_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11622_ (.A1(_03643_),
    .A2(_02024_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11623_ (.A1(\channels.pw3[4] ),
    .A2(_03727_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11624_ (.I(_03717_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11625_ (.A1(_03647_),
    .A2(_03729_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11626_ (.A1(_03728_),
    .A2(_03730_),
    .B(_03652_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11627_ (.A1(\channels.pw3[5] ),
    .A2(_03718_),
    .B(_03723_),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11628_ (.A1(_03693_),
    .A2(_03729_),
    .B(_03731_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11629_ (.I(_03722_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11630_ (.A1(\channels.pw3[6] ),
    .A2(_03718_),
    .B(_03732_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11631_ (.A1(_03695_),
    .A2(_03729_),
    .B(_03733_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11632_ (.A1(\channels.pw3[7] ),
    .A2(_03718_),
    .B(_03732_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11633_ (.A1(_03697_),
    .A2(_03729_),
    .B(_03734_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11634_ (.I(_01750_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11635_ (.A1(_03658_),
    .A2(_01856_),
    .Z(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11636_ (.I(_03736_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11637_ (.I(_03737_),
    .Z(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11638_ (.I(_03736_),
    .Z(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11639_ (.A1(\channels.pw2[0] ),
    .A2(_03739_),
    .B(_03732_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11640_ (.A1(_03735_),
    .A2(_03738_),
    .B(_03740_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11641_ (.A1(\channels.pw2[1] ),
    .A2(_03739_),
    .B(_03732_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11642_ (.A1(_03683_),
    .A2(_03738_),
    .B(_03741_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11643_ (.I(_03722_),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11644_ (.A1(\channels.pw2[2] ),
    .A2(_03739_),
    .B(_03742_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11645_ (.A1(_03685_),
    .A2(_03738_),
    .B(_03743_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11646_ (.A1(\channels.pw2[3] ),
    .A2(_03739_),
    .B(_03742_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11647_ (.A1(_03707_),
    .A2(_03738_),
    .B(_03744_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11648_ (.A1(_02352_),
    .A2(_02008_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11649_ (.A1(\channels.pw2[4] ),
    .A2(_03745_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11650_ (.I(_03646_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11651_ (.I(_03736_),
    .Z(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11652_ (.A1(_03747_),
    .A2(_03748_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11653_ (.I(_03651_),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11654_ (.A1(_03746_),
    .A2(_03749_),
    .B(_03750_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11655_ (.A1(\channels.pw2[5] ),
    .A2(_03737_),
    .B(_03742_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11656_ (.A1(_03693_),
    .A2(_03748_),
    .B(_03751_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11657_ (.A1(\channels.pw2[6] ),
    .A2(_03737_),
    .B(_03742_),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11658_ (.A1(_03695_),
    .A2(_03748_),
    .B(_03752_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11659_ (.I(_03722_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11660_ (.A1(\channels.pw2[7] ),
    .A2(_03737_),
    .B(_03753_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11661_ (.A1(_03697_),
    .A2(_03748_),
    .B(_03754_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11662_ (.A1(_01103_),
    .A2(_03497_),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11663_ (.I(_03755_),
    .Z(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11664_ (.I(_01079_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11665_ (.I(_03757_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11666_ (.I(_03758_),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11667_ (.I(_03759_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11668_ (.I(_01761_),
    .Z(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11669_ (.I(_03761_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11670_ (.A1(\channels.clk_div[0] ),
    .A2(_03760_),
    .B(_03762_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11671_ (.A1(_03756_),
    .A2(_03763_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11672_ (.I(_01274_),
    .Z(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11673_ (.A1(_03764_),
    .A2(_03756_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11674_ (.I(_01760_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11675_ (.I(_03766_),
    .Z(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11676_ (.A1(_03764_),
    .A2(_03755_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11677_ (.A1(_03767_),
    .A2(_03768_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11678_ (.A1(_03765_),
    .A2(_03769_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11679_ (.A1(_01593_),
    .A2(_03768_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11680_ (.A1(_01945_),
    .A2(_03770_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11681_ (.I(_02841_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11682_ (.I(_03771_),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11683_ (.I(_01329_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11684_ (.I(_03133_),
    .Z(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11685_ (.I(_03041_),
    .Z(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11686_ (.I(_02723_),
    .Z(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11687_ (.I(_02689_),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11688_ (.A1(_03777_),
    .A2(_03771_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11689_ (.A1(_03776_),
    .A2(_03778_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11690_ (.A1(_03775_),
    .A2(_03779_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11691_ (.A1(_03098_),
    .A2(_03549_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11692_ (.I(_03781_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11693_ (.A1(_03544_),
    .A2(_03780_),
    .A3(_03782_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11694_ (.A1(_03774_),
    .A2(_03783_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11695_ (.A1(_03539_),
    .A2(_03540_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11696_ (.I(_03785_),
    .Z(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11697_ (.A1(\channels.sus_rel1[5] ),
    .A2(_01304_),
    .Z(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11698_ (.A1(\channels.sus_rel3[5] ),
    .A2(_01092_),
    .B1(_01291_),
    .B2(\channels.sus_rel2[5] ),
    .C(_03787_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11699_ (.A1(_03549_),
    .A2(_03788_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11700_ (.A1(_03777_),
    .A2(_03788_),
    .B(_03789_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11701_ (.A1(\channels.sus_rel1[4] ),
    .A2(_01304_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11702_ (.A1(\channels.sus_rel3[4] ),
    .A2(_01092_),
    .B1(_01291_),
    .B2(\channels.sus_rel2[4] ),
    .C(_03791_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11703_ (.I0(_02713_),
    .I1(_03548_),
    .S(_03792_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11704_ (.A1(\channels.sus_rel3[7] ),
    .A2(_01091_),
    .Z(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11705_ (.A1(\channels.sus_rel2[7] ),
    .A2(_01291_),
    .B1(_01305_),
    .B2(\channels.sus_rel1[7] ),
    .C(_03794_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11706_ (.A1(_01178_),
    .A2(_02534_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _11707_ (.A1(_01178_),
    .A2(_02535_),
    .B(_03796_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11708_ (.A1(\channels.sus_rel3[6] ),
    .A2(_01092_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11709_ (.A1(\channels.sus_rel2[6] ),
    .A2(_01290_),
    .B1(_01304_),
    .B2(\channels.sus_rel1[6] ),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _11710_ (.A1(_03798_),
    .A2(_03799_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11711_ (.A1(_03797_),
    .A2(_03090_),
    .B1(_03800_),
    .B2(_03776_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _11712_ (.A1(_03548_),
    .A2(_02713_),
    .B1(_03133_),
    .B2(_03795_),
    .C(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11713_ (.A1(_03777_),
    .A2(_02754_),
    .B1(_03795_),
    .B2(_03041_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11714_ (.A1(_03545_),
    .A2(_03544_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11715_ (.A1(_03544_),
    .A2(_03800_),
    .B(_03803_),
    .C(_03804_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11716_ (.A1(_03790_),
    .A2(_03793_),
    .A3(_03802_),
    .A4(_03805_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11717_ (.A1(_03559_),
    .A2(_03784_),
    .B1(_03786_),
    .B2(_03806_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11718_ (.A1(_03543_),
    .A2(_03807_),
    .Z(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11719_ (.I(_01435_),
    .Z(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11720_ (.A1(\channels.sus_rel3[0] ),
    .A2(_01449_),
    .B1(_03809_),
    .B2(\channels.sus_rel2[0] ),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11721_ (.I(_01407_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11722_ (.I(_01287_),
    .Z(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11723_ (.I(_03785_),
    .Z(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11724_ (.I(_03813_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11725_ (.A1(\channels.atk_dec3[0] ),
    .A2(_03811_),
    .B1(_03812_),
    .B2(\channels.atk_dec2[0] ),
    .C(_03814_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11726_ (.A1(_03786_),
    .A2(_03810_),
    .B(_03815_),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11727_ (.I(_01300_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11728_ (.I0(\channels.atk_dec1[0] ),
    .I1(\channels.sus_rel1[0] ),
    .S(_03813_),
    .Z(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11729_ (.A1(_03817_),
    .A2(_03818_),
    .Z(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11730_ (.I(_03541_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11731_ (.A1(\channels.atk_dec3[4] ),
    .A2(_01089_),
    .B1(_03809_),
    .B2(\channels.atk_dec2[4] ),
    .C1(_01301_),
    .C2(\channels.atk_dec1[4] ),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11732_ (.A1(_03820_),
    .A2(_03821_),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _11733_ (.A1(_03542_),
    .A2(_03816_),
    .A3(_03819_),
    .B(_03822_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11734_ (.A1(\channels.atk_dec3[1] ),
    .A2(_01088_),
    .B1(_01435_),
    .B2(\channels.atk_dec2[1] ),
    .ZN(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11735_ (.A1(\channels.sus_rel3[1] ),
    .A2(_01088_),
    .B1(_01435_),
    .B2(\channels.sus_rel2[1] ),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11736_ (.I0(_03824_),
    .I1(_03825_),
    .S(_03814_),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11737_ (.I0(\channels.atk_dec1[1] ),
    .I1(\channels.sus_rel1[1] ),
    .S(_03813_),
    .Z(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11738_ (.A1(_03817_),
    .A2(_03827_),
    .B(_03541_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _11739_ (.A1(\channels.atk_dec3[5] ),
    .A2(_01089_),
    .B1(_03809_),
    .B2(\channels.atk_dec2[5] ),
    .C1(_01301_),
    .C2(\channels.atk_dec1[5] ),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _11740_ (.A1(_03826_),
    .A2(_03828_),
    .B1(_03829_),
    .B2(_03820_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11741_ (.I(_03830_),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11742_ (.I(_03831_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11743_ (.A1(_03823_),
    .A2(_03832_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11744_ (.I(_03823_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11745_ (.A1(\channels.sus_rel3[2] ),
    .A2(_03811_),
    .B1(_01288_),
    .B2(\channels.sus_rel2[2] ),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11746_ (.A1(\channels.atk_dec3[2] ),
    .A2(_03811_),
    .B1(_01288_),
    .B2(\channels.atk_dec2[2] ),
    .C(_03814_),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11747_ (.A1(_03786_),
    .A2(_03835_),
    .B(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11748_ (.I0(\channels.atk_dec1[2] ),
    .I1(\channels.sus_rel1[2] ),
    .S(_03813_),
    .Z(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11749_ (.A1(_03817_),
    .A2(_03838_),
    .Z(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11750_ (.A1(\channels.atk_dec3[6] ),
    .A2(_01449_),
    .B1(_03812_),
    .B2(\channels.atk_dec2[6] ),
    .C1(_01301_),
    .C2(\channels.atk_dec1[6] ),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11751_ (.A1(_03820_),
    .A2(_03840_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _11752_ (.A1(_03542_),
    .A2(_03837_),
    .A3(_03839_),
    .B(_03841_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11753_ (.I(_03842_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11754_ (.A1(_03834_),
    .A2(_03843_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11755_ (.A1(_03832_),
    .A2(_03844_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11756_ (.A1(\channels.atk_dec3[3] ),
    .A2(_01449_),
    .B1(_03812_),
    .B2(\channels.atk_dec2[3] ),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11757_ (.A1(\channels.sus_rel3[3] ),
    .A2(_03811_),
    .B1(_03812_),
    .B2(\channels.sus_rel2[3] ),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11758_ (.I0(_03846_),
    .I1(_03847_),
    .S(_03786_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11759_ (.I0(\channels.atk_dec1[3] ),
    .I1(\channels.sus_rel1[3] ),
    .S(_03814_),
    .Z(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11760_ (.A1(_01302_),
    .A2(_03849_),
    .B(_03820_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11761_ (.A1(\channels.atk_dec3[7] ),
    .A2(_01089_),
    .B1(_03809_),
    .B2(\channels.atk_dec2[7] ),
    .C1(_03817_),
    .C2(\channels.atk_dec1[7] ),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11762_ (.A1(_03848_),
    .A2(_03850_),
    .B1(_03851_),
    .B2(_03542_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11763_ (.I(_03852_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11764_ (.A1(_03843_),
    .A2(_03853_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11765_ (.A1(_03842_),
    .A2(_03852_),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11766_ (.A1(_03854_),
    .A2(_03855_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11767_ (.A1(_03830_),
    .A2(_03843_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11768_ (.A1(_03845_),
    .A2(_03856_),
    .B(_03857_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11769_ (.A1(_03833_),
    .A2(_03858_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11770_ (.I(_01160_),
    .Z(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11771_ (.I(_03860_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11772_ (.I0(\channels.env_counter[0][2] ),
    .I1(\channels.env_counter[1][2] ),
    .I2(\channels.env_counter[2][2] ),
    .I3(\channels.env_counter[3][2] ),
    .S0(_03861_),
    .S1(_01181_),
    .Z(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _11773_ (.A1(_03859_),
    .A2(_03862_),
    .Z(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11774_ (.I(_03852_),
    .Z(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11775_ (.I(_03864_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11776_ (.I(_03823_),
    .Z(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11777_ (.A1(_03831_),
    .A2(_03842_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11778_ (.A1(_03857_),
    .A2(_03867_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11779_ (.A1(_03866_),
    .A2(_03868_),
    .Z(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11780_ (.A1(_03865_),
    .A2(_03869_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11781_ (.I(_01176_),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11782_ (.I0(\channels.env_counter[0][9] ),
    .I1(\channels.env_counter[1][9] ),
    .I2(\channels.env_counter[2][9] ),
    .I3(\channels.env_counter[3][9] ),
    .S0(_03861_),
    .S1(_03871_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11783_ (.A1(_03870_),
    .A2(_03872_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11784_ (.I(_03842_),
    .Z(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11785_ (.A1(_03874_),
    .A2(_03864_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11786_ (.A1(_03834_),
    .A2(_03864_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11787_ (.A1(_03875_),
    .A2(_03876_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11788_ (.I(_03877_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11789_ (.I(_03830_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11790_ (.A1(_03866_),
    .A2(_03879_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11791_ (.A1(_03866_),
    .A2(_03868_),
    .B(_03853_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11792_ (.A1(_03878_),
    .A2(_03880_),
    .B(_03881_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11793_ (.I0(\channels.env_counter[0][6] ),
    .I1(\channels.env_counter[1][6] ),
    .I2(\channels.env_counter[2][6] ),
    .I3(\channels.env_counter[3][6] ),
    .S0(_03861_),
    .S1(_03871_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11794_ (.A1(_03882_),
    .A2(_03883_),
    .Z(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11795_ (.A1(_03863_),
    .A2(_03873_),
    .A3(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11796_ (.I(_03844_),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11797_ (.I(_03886_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11798_ (.A1(_03866_),
    .A2(_03856_),
    .B(_03887_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11799_ (.A1(_03879_),
    .A2(_03888_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11800_ (.I0(\channels.env_counter[0][5] ),
    .I1(\channels.env_counter[1][5] ),
    .I2(\channels.env_counter[2][5] ),
    .I3(\channels.env_counter[3][5] ),
    .S0(_01162_),
    .S1(_01181_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11801_ (.I(_03890_),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11802_ (.A1(_03889_),
    .A2(_03891_),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11803_ (.A1(_03879_),
    .A2(_03874_),
    .B(_03834_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11804_ (.A1(_03865_),
    .A2(_03868_),
    .B(_03893_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11805_ (.I0(\channels.env_counter[0][4] ),
    .I1(\channels.env_counter[1][4] ),
    .I2(\channels.env_counter[2][4] ),
    .I3(\channels.env_counter[3][4] ),
    .S0(_03860_),
    .S1(_01177_),
    .Z(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _11806_ (.A1(_03894_),
    .A2(_03895_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11807_ (.A1(_03823_),
    .A2(_03874_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11808_ (.A1(_03830_),
    .A2(_03897_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11809_ (.A1(_03833_),
    .A2(_03898_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11810_ (.A1(_03853_),
    .A2(_03899_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11811_ (.A1(_03833_),
    .A2(_03854_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11812_ (.A1(_03900_),
    .A2(_03901_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11813_ (.I0(\channels.env_counter[0][1] ),
    .I1(\channels.env_counter[1][1] ),
    .I2(\channels.env_counter[2][1] ),
    .I3(\channels.env_counter[3][1] ),
    .S0(_03860_),
    .S1(_01177_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11814_ (.A1(_03902_),
    .A2(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11815_ (.A1(_03892_),
    .A2(_03896_),
    .A3(_03904_),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11816_ (.A1(_03832_),
    .A2(_03887_),
    .B(_03897_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11817_ (.A1(_03875_),
    .A2(_03880_),
    .B1(_03906_),
    .B2(_03865_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _11818_ (.I0(\channels.env_counter[0][0] ),
    .I1(\channels.env_counter[1][0] ),
    .I2(\channels.env_counter[2][0] ),
    .I3(\channels.env_counter[3][0] ),
    .S0(_01161_),
    .S1(_01177_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11819_ (.I(_03908_),
    .Z(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11820_ (.A1(_03907_),
    .A2(_03909_),
    .Z(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11821_ (.A1(_03907_),
    .A2(_03909_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11822_ (.A1(_03902_),
    .A2(_03903_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11823_ (.I(_03877_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11824_ (.A1(_03833_),
    .A2(_03874_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11825_ (.I(_01159_),
    .Z(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _11826_ (.I0(\channels.env_counter[0][3] ),
    .I1(\channels.env_counter[1][3] ),
    .I2(\channels.env_counter[2][3] ),
    .I3(\channels.env_counter[3][3] ),
    .S0(_03915_),
    .S1(_01176_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11827_ (.I(_03916_),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11828_ (.A1(_03913_),
    .A2(_03914_),
    .B(_03917_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11829_ (.I(_03864_),
    .Z(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11830_ (.A1(_03919_),
    .A2(_03898_),
    .A3(_03867_),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11831_ (.I0(\channels.env_counter[0][10] ),
    .I1(\channels.env_counter[1][10] ),
    .I2(\channels.env_counter[2][10] ),
    .I3(\channels.env_counter[3][10] ),
    .S0(_03915_),
    .S1(_01180_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11832_ (.A1(_03913_),
    .A2(_03914_),
    .A3(_03916_),
    .B1(_03920_),
    .B2(_03921_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11833_ (.I(_03922_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11834_ (.A1(_03889_),
    .A2(_03890_),
    .B(_03918_),
    .C(_03923_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _11835_ (.A1(_03910_),
    .A2(_03911_),
    .A3(_03912_),
    .A4(_03924_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11836_ (.A1(_03919_),
    .A2(_03867_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _11837_ (.I0(\channels.env_counter[0][11] ),
    .I1(\channels.env_counter[1][11] ),
    .I2(\channels.env_counter[2][11] ),
    .I3(\channels.env_counter[3][11] ),
    .S0(_01160_),
    .S1(_01175_),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11838_ (.A1(_03886_),
    .A2(_03926_),
    .A3(_03927_),
    .Z(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11839_ (.I(_03927_),
    .Z(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11840_ (.A1(_03886_),
    .A2(_03926_),
    .B(_03929_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _11841_ (.A1(_03832_),
    .A2(_03886_),
    .B1(_03855_),
    .B2(_03913_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11842_ (.I0(\channels.env_counter[0][7] ),
    .I1(\channels.env_counter[1][7] ),
    .I2(\channels.env_counter[2][7] ),
    .I3(\channels.env_counter[3][7] ),
    .S0(_01161_),
    .S1(_03871_),
    .Z(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11843_ (.A1(_03931_),
    .A2(_03932_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11844_ (.I0(\channels.env_counter[0][8] ),
    .I1(\channels.env_counter[1][8] ),
    .I2(\channels.env_counter[2][8] ),
    .I3(\channels.env_counter[3][8] ),
    .S0(_03861_),
    .S1(_01181_),
    .Z(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11845_ (.I(_03857_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11846_ (.I0(_03935_),
    .I1(_03845_),
    .S(_03865_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11847_ (.A1(_03934_),
    .A2(_03936_),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _11848_ (.I0(\channels.env_counter[0][12] ),
    .I1(\channels.env_counter[1][12] ),
    .I2(\channels.env_counter[2][12] ),
    .I3(\channels.env_counter[3][12] ),
    .S0(_01160_),
    .S1(_01176_),
    .Z(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11849_ (.A1(_03935_),
    .A2(_03876_),
    .B(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11850_ (.I(_03938_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11851_ (.A1(_03935_),
    .A2(_03876_),
    .A3(_03940_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11852_ (.A1(_03933_),
    .A2(_03937_),
    .A3(_03939_),
    .A4(_03941_),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11853_ (.I(_03934_),
    .Z(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11854_ (.A1(_03919_),
    .A2(_03897_),
    .Z(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11855_ (.I0(\channels.env_counter[0][13] ),
    .I1(\channels.env_counter[1][13] ),
    .S(_03915_),
    .Z(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11856_ (.I(\channels.env_counter[2][13] ),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11857_ (.A1(_03860_),
    .A2(\channels.env_counter[3][13] ),
    .ZN(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11858_ (.A1(_01161_),
    .A2(_03946_),
    .B(_03947_),
    .C(_01180_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11859_ (.A1(_03871_),
    .A2(_03945_),
    .B(_03948_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11860_ (.A1(_03944_),
    .A2(_03949_),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11861_ (.A1(_03920_),
    .A2(_03921_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11862_ (.A1(_03944_),
    .A2(_03949_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11863_ (.A1(_03879_),
    .A2(_03843_),
    .A3(_03919_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _11864_ (.I0(\channels.env_counter[0][14] ),
    .I1(\channels.env_counter[1][14] ),
    .I2(\channels.env_counter[2][14] ),
    .I3(\channels.env_counter[3][14] ),
    .S0(_03915_),
    .S1(_01180_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11865_ (.A1(_03953_),
    .A2(_03954_),
    .Z(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11866_ (.A1(_03953_),
    .A2(_03954_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11867_ (.A1(_03952_),
    .A2(_03955_),
    .A3(_03956_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11868_ (.A1(_01594_),
    .A2(_03950_),
    .A3(_03951_),
    .A4(_03957_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11869_ (.A1(_03931_),
    .A2(_03932_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11870_ (.I(_03959_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11871_ (.A1(_03943_),
    .A2(_03936_),
    .B(_03958_),
    .C(_03960_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11872_ (.A1(_03928_),
    .A2(_03930_),
    .A3(_03942_),
    .A4(_03961_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11873_ (.A1(_03885_),
    .A2(_03905_),
    .A3(_03925_),
    .A4(_03962_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11874_ (.I(_03963_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11875_ (.A1(_03808_),
    .A2(_03964_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11876_ (.I(_03965_),
    .Z(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11877_ (.A1(_03773_),
    .A2(_03966_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11878_ (.I(_03967_),
    .Z(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11879_ (.A1(_03773_),
    .A2(_03966_),
    .B(_03650_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11880_ (.I(_03969_),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11881_ (.A1(\channels.env_vol[0][0] ),
    .A2(_03970_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11882_ (.A1(_03772_),
    .A2(_03968_),
    .B(_03971_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11883_ (.A1(_03546_),
    .A2(_03778_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11884_ (.A1(_03807_),
    .A2(_03963_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11885_ (.I(_03973_),
    .Z(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11886_ (.I(_03974_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11887_ (.A1(_03972_),
    .A2(_03975_),
    .Z(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11888_ (.A1(\channels.env_vol[0][1] ),
    .A2(_03970_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11889_ (.A1(_03968_),
    .A2(_03976_),
    .B(_03977_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11890_ (.A1(_03777_),
    .A2(_03772_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11891_ (.I(_03973_),
    .Z(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11892_ (.A1(_03778_),
    .A2(_03974_),
    .ZN(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11893_ (.A1(_03978_),
    .A2(_03979_),
    .B(_03980_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11894_ (.A1(_03776_),
    .A2(_03981_),
    .Z(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11895_ (.A1(\channels.env_vol[0][2] ),
    .A2(_03970_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11896_ (.A1(_03968_),
    .A2(_03982_),
    .B(_03983_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11897_ (.A1(_03545_),
    .A2(_03979_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11898_ (.A1(_03978_),
    .A2(_03979_),
    .B1(_03984_),
    .B2(_03779_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11899_ (.A1(_03797_),
    .A2(_03985_),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11900_ (.A1(\channels.env_vol[0][3] ),
    .A2(_03970_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11901_ (.A1(_03968_),
    .A2(_03986_),
    .B(_03987_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11902_ (.I(_03967_),
    .Z(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11903_ (.I(_03780_),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11904_ (.A1(_03547_),
    .A2(_03979_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11905_ (.A1(_03989_),
    .A2(_03975_),
    .B(_03990_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11906_ (.A1(_03548_),
    .A2(_03991_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11907_ (.I(_03969_),
    .Z(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11908_ (.A1(\channels.env_vol[0][4] ),
    .A2(_03993_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11909_ (.A1(_03988_),
    .A2(_03992_),
    .B(_03994_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11910_ (.A1(_03551_),
    .A2(_03781_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11911_ (.A1(_02754_),
    .A2(_03547_),
    .B(_03995_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11912_ (.I(_03989_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11913_ (.A1(_03549_),
    .A2(_03997_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11914_ (.A1(_03550_),
    .A2(_03781_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11915_ (.A1(_03989_),
    .A2(_03999_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11916_ (.A1(_03998_),
    .A2(_04000_),
    .B(_03975_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11917_ (.A1(_03975_),
    .A2(_03996_),
    .B(_04001_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11918_ (.A1(\channels.env_vol[0][5] ),
    .A2(_03993_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11919_ (.A1(_03988_),
    .A2(_04002_),
    .B(_04003_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11920_ (.A1(_03989_),
    .A2(_03782_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11921_ (.I0(_04004_),
    .I1(_03551_),
    .S(_03974_),
    .Z(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11922_ (.A1(_03130_),
    .A2(_04005_),
    .Z(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11923_ (.A1(\channels.env_vol[0][6] ),
    .A2(_03993_),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11924_ (.A1(_03988_),
    .A2(_04006_),
    .B(_04007_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11925_ (.I0(_03783_),
    .I1(_03552_),
    .S(_03974_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11926_ (.A1(_03774_),
    .A2(_04008_),
    .Z(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11927_ (.A1(\channels.env_vol[0][7] ),
    .A2(_03993_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11928_ (.A1(_03988_),
    .A2(_04009_),
    .B(_04010_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11929_ (.A1(_03907_),
    .A2(_03908_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11930_ (.A1(_03952_),
    .A2(_03955_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11931_ (.A1(_04011_),
    .A2(_03950_),
    .A3(_04012_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11932_ (.A1(_03934_),
    .A2(_03936_),
    .B(_04013_),
    .C(_03911_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11933_ (.A1(_03959_),
    .A2(_03933_),
    .A3(_03937_),
    .A4(_04014_),
    .Z(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11934_ (.A1(_03889_),
    .A2(_03890_),
    .B(_03912_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11935_ (.A1(_03889_),
    .A2(_03891_),
    .B(_04016_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11936_ (.A1(_03873_),
    .A2(_03896_),
    .A3(_03904_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11937_ (.A1(_03920_),
    .A2(_03921_),
    .B(_03928_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11938_ (.I(_04019_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11939_ (.A1(_03913_),
    .A2(_03914_),
    .A3(_03917_),
    .Z(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11940_ (.A1(_03930_),
    .A2(_03951_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11941_ (.A1(_01594_),
    .A2(_03939_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11942_ (.A1(_03935_),
    .A2(_03876_),
    .A3(_03940_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _11943_ (.A1(_04022_),
    .A2(_04023_),
    .A3(_04024_),
    .A4(_03956_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11944_ (.A1(_04020_),
    .A2(_03918_),
    .A3(_04021_),
    .A4(_04025_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11945_ (.A1(_03884_),
    .A2(_04026_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11946_ (.A1(_04017_),
    .A2(_04018_),
    .A3(_04027_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _11947_ (.A1(_03863_),
    .A2(_04015_),
    .A3(_04028_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11948_ (.A1(_01195_),
    .A2(_01201_),
    .A3(_01208_),
    .A4(_01233_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11949_ (.A1(_03543_),
    .A2(_04030_),
    .B(_01595_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11950_ (.A1(_04029_),
    .A2(_04031_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11951_ (.I(_04032_),
    .Z(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11952_ (.A1(_02358_),
    .A2(_04033_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11953_ (.I(_04034_),
    .Z(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11954_ (.I(_04035_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11955_ (.I(_03964_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11956_ (.A1(_03909_),
    .A2(_04037_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11957_ (.A1(_01591_),
    .A2(_04033_),
    .B(_01825_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11958_ (.I(_04039_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11959_ (.I(_04040_),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11960_ (.A1(\channels.env_counter[2][0] ),
    .A2(_04041_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11961_ (.A1(_04036_),
    .A2(_04038_),
    .B(_04042_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11962_ (.A1(_03908_),
    .A2(_03903_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11963_ (.A1(_03909_),
    .A2(_03903_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11964_ (.A1(_04037_),
    .A2(_04043_),
    .A3(_04044_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11965_ (.A1(\channels.env_counter[2][1] ),
    .A2(_04041_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11966_ (.A1(_04036_),
    .A2(_04045_),
    .B(_04046_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11967_ (.I(_04029_),
    .Z(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11968_ (.A1(_03862_),
    .A2(_04043_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11969_ (.A1(_04047_),
    .A2(_04048_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11970_ (.A1(\channels.env_counter[2][2] ),
    .A2(_04041_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11971_ (.A1(_04036_),
    .A2(_04049_),
    .B(_04050_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11972_ (.A1(_03862_),
    .A2(_03917_),
    .A3(_04043_),
    .Z(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11973_ (.A1(_03862_),
    .A2(_04043_),
    .B(_03917_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11974_ (.A1(_04037_),
    .A2(_04051_),
    .A3(_04052_),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11975_ (.A1(\channels.env_counter[2][3] ),
    .A2(_04041_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11976_ (.A1(_04036_),
    .A2(_04053_),
    .B(_04054_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11977_ (.I(_04034_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11978_ (.A1(_03895_),
    .A2(_04051_),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11979_ (.A1(_04047_),
    .A2(_04056_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11980_ (.I(_04039_),
    .Z(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11981_ (.A1(\channels.env_counter[2][4] ),
    .A2(_04058_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11982_ (.A1(_04055_),
    .A2(_04057_),
    .B(_04059_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11983_ (.A1(_03891_),
    .A2(_03895_),
    .A3(_04051_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11984_ (.A1(_03895_),
    .A2(_04051_),
    .B(_03891_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11985_ (.A1(_04037_),
    .A2(_04060_),
    .A3(_04061_),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11986_ (.A1(\channels.env_counter[2][5] ),
    .A2(_04058_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11987_ (.A1(_04055_),
    .A2(_04062_),
    .B(_04063_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11988_ (.A1(_03883_),
    .A2(_04060_),
    .Z(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11989_ (.A1(_04047_),
    .A2(_04064_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11990_ (.A1(\channels.env_counter[2][6] ),
    .A2(_04058_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11991_ (.A1(_04055_),
    .A2(_04065_),
    .B(_04066_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11992_ (.A1(_03932_),
    .A2(_03883_),
    .A3(_04060_),
    .Z(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11993_ (.A1(_03883_),
    .A2(_04060_),
    .B(_03932_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _11994_ (.A1(_03964_),
    .A2(_04067_),
    .A3(_04068_),
    .Z(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11995_ (.A1(\channels.env_counter[2][7] ),
    .A2(_04058_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11996_ (.A1(_04055_),
    .A2(_04069_),
    .B(_04070_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11997_ (.I(_04034_),
    .Z(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11998_ (.I(_04029_),
    .Z(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11999_ (.A1(_03943_),
    .A2(_04067_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12000_ (.A1(_03943_),
    .A2(_04067_),
    .Z(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12001_ (.A1(_04072_),
    .A2(_04073_),
    .A3(_04074_),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12002_ (.I(_04039_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12003_ (.A1(\channels.env_counter[2][8] ),
    .A2(_04076_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12004_ (.A1(_04071_),
    .A2(_04075_),
    .B(_04077_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12005_ (.A1(_03872_),
    .A2(_04073_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12006_ (.A1(_04047_),
    .A2(_04078_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12007_ (.A1(\channels.env_counter[2][9] ),
    .A2(_04076_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12008_ (.A1(_04071_),
    .A2(_04079_),
    .B(_04080_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12009_ (.I(_03921_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12010_ (.A1(_03943_),
    .A2(_03872_),
    .A3(_04067_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12011_ (.A1(_04081_),
    .A2(_04082_),
    .Z(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12012_ (.A1(_04072_),
    .A2(_04083_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12013_ (.A1(\channels.env_counter[2][10] ),
    .A2(_04076_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12014_ (.A1(_04071_),
    .A2(_04084_),
    .B(_04085_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12015_ (.A1(_04081_),
    .A2(_04082_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12016_ (.A1(_03929_),
    .A2(_04086_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12017_ (.A1(_03929_),
    .A2(_04086_),
    .Z(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12018_ (.A1(_04029_),
    .A2(_04087_),
    .A3(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12019_ (.A1(\channels.env_counter[2][11] ),
    .A2(_04076_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12020_ (.A1(_04071_),
    .A2(_04089_),
    .B(_04090_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12021_ (.A1(_03940_),
    .A2(_04087_),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12022_ (.A1(_04072_),
    .A2(_04091_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12023_ (.A1(\channels.env_counter[2][12] ),
    .A2(_04040_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12024_ (.A1(_04035_),
    .A2(_04092_),
    .B(_04093_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12025_ (.A1(_03929_),
    .A2(_03940_),
    .A3(_04086_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12026_ (.A1(_03949_),
    .A2(_04094_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12027_ (.A1(_04072_),
    .A2(_04095_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12028_ (.A1(\channels.env_counter[2][13] ),
    .A2(_04040_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12029_ (.A1(_04035_),
    .A2(_04096_),
    .B(_04097_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12030_ (.A1(_03949_),
    .A2(_04094_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12031_ (.A1(_03954_),
    .A2(_04098_),
    .B(_03964_),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12032_ (.A1(_03954_),
    .A2(_04098_),
    .B(_04099_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12033_ (.A1(\channels.env_counter[2][14] ),
    .A2(_04040_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12034_ (.A1(_04035_),
    .A2(_04100_),
    .B(_04101_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12035_ (.A1(_02365_),
    .A2(_04033_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12036_ (.I(_04102_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12037_ (.I(_04103_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12038_ (.A1(_03764_),
    .A2(_04032_),
    .B(_01825_),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12039_ (.I(_04105_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12040_ (.I(_04106_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12041_ (.A1(\channels.env_counter[1][0] ),
    .A2(_04107_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12042_ (.A1(_04038_),
    .A2(_04104_),
    .B(_04108_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12043_ (.A1(\channels.env_counter[1][1] ),
    .A2(_04107_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12044_ (.A1(_04045_),
    .A2(_04104_),
    .B(_04109_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12045_ (.A1(\channels.env_counter[1][2] ),
    .A2(_04107_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12046_ (.A1(_04049_),
    .A2(_04104_),
    .B(_04110_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12047_ (.A1(\channels.env_counter[1][3] ),
    .A2(_04107_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12048_ (.A1(_04053_),
    .A2(_04104_),
    .B(_04111_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12049_ (.I(_04102_),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12050_ (.I(_04105_),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12051_ (.A1(\channels.env_counter[1][4] ),
    .A2(_04113_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12052_ (.A1(_04057_),
    .A2(_04112_),
    .B(_04114_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12053_ (.A1(\channels.env_counter[1][5] ),
    .A2(_04113_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12054_ (.A1(_04062_),
    .A2(_04112_),
    .B(_04115_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12055_ (.A1(\channels.env_counter[1][6] ),
    .A2(_04113_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12056_ (.A1(_04065_),
    .A2(_04112_),
    .B(_04116_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12057_ (.A1(\channels.env_counter[1][7] ),
    .A2(_04113_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12058_ (.A1(_04069_),
    .A2(_04112_),
    .B(_04117_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12059_ (.I(_04102_),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12060_ (.I(_04105_),
    .Z(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12061_ (.A1(\channels.env_counter[1][8] ),
    .A2(_04119_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12062_ (.A1(_04075_),
    .A2(_04118_),
    .B(_04120_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12063_ (.A1(\channels.env_counter[1][9] ),
    .A2(_04119_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12064_ (.A1(_04079_),
    .A2(_04118_),
    .B(_04121_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12065_ (.A1(\channels.env_counter[1][10] ),
    .A2(_04119_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12066_ (.A1(_04084_),
    .A2(_04118_),
    .B(_04122_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12067_ (.A1(\channels.env_counter[1][11] ),
    .A2(_04119_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12068_ (.A1(_04089_),
    .A2(_04118_),
    .B(_04123_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12069_ (.A1(\channels.env_counter[1][12] ),
    .A2(_04106_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12070_ (.A1(_04092_),
    .A2(_04103_),
    .B(_04124_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12071_ (.A1(\channels.env_counter[1][13] ),
    .A2(_04106_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12072_ (.A1(_04096_),
    .A2(_04103_),
    .B(_04125_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12073_ (.A1(\channels.env_counter[1][14] ),
    .A2(_04106_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12074_ (.A1(_04100_),
    .A2(_04103_),
    .B(_04126_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12075_ (.I(\channels.adsr_state[3][0] ),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12076_ (.I(_04127_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12077_ (.I(\channels.adsr_state[3][1] ),
    .Z(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12078_ (.I(_04128_),
    .Z(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _12079_ (.A1(\clk_ctr[0] ),
    .A2(_02356_),
    .A3(_03760_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12080_ (.I(_03561_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12081_ (.A1(_01072_),
    .A2(\clk_ctr[1] ),
    .Z(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _12082_ (.A1(_04129_),
    .A2(_03760_),
    .A3(_04130_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12083_ (.A1(_03773_),
    .A2(_04033_),
    .ZN(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12084_ (.I(_04131_),
    .Z(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12085_ (.I(_04132_),
    .Z(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12086_ (.A1(_01329_),
    .A2(_04032_),
    .B(_01825_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12087_ (.I(_04134_),
    .Z(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12088_ (.I(_04135_),
    .Z(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12089_ (.A1(\channels.env_counter[0][0] ),
    .A2(_04136_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12090_ (.A1(_04038_),
    .A2(_04133_),
    .B(_04137_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12091_ (.A1(\channels.env_counter[0][1] ),
    .A2(_04136_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12092_ (.A1(_04045_),
    .A2(_04133_),
    .B(_04138_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12093_ (.A1(\channels.env_counter[0][2] ),
    .A2(_04136_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12094_ (.A1(_04049_),
    .A2(_04133_),
    .B(_04139_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12095_ (.A1(\channels.env_counter[0][3] ),
    .A2(_04136_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12096_ (.A1(_04053_),
    .A2(_04133_),
    .B(_04140_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12097_ (.I(_04131_),
    .Z(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12098_ (.I(_04134_),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12099_ (.A1(\channels.env_counter[0][4] ),
    .A2(_04142_),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12100_ (.A1(_04057_),
    .A2(_04141_),
    .B(_04143_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12101_ (.A1(\channels.env_counter[0][5] ),
    .A2(_04142_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12102_ (.A1(_04062_),
    .A2(_04141_),
    .B(_04144_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12103_ (.A1(\channels.env_counter[0][6] ),
    .A2(_04142_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12104_ (.A1(_04065_),
    .A2(_04141_),
    .B(_04145_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12105_ (.A1(\channels.env_counter[0][7] ),
    .A2(_04142_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12106_ (.A1(_04069_),
    .A2(_04141_),
    .B(_04146_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12107_ (.I(_04131_),
    .Z(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12108_ (.I(_04134_),
    .Z(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12109_ (.A1(\channels.env_counter[0][8] ),
    .A2(_04148_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12110_ (.A1(_04075_),
    .A2(_04147_),
    .B(_04149_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12111_ (.A1(\channels.env_counter[0][9] ),
    .A2(_04148_),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12112_ (.A1(_04079_),
    .A2(_04147_),
    .B(_04150_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12113_ (.A1(\channels.env_counter[0][10] ),
    .A2(_04148_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12114_ (.A1(_04084_),
    .A2(_04147_),
    .B(_04151_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12115_ (.A1(\channels.env_counter[0][11] ),
    .A2(_04148_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12116_ (.A1(_04089_),
    .A2(_04147_),
    .B(_04152_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12117_ (.A1(\channels.env_counter[0][12] ),
    .A2(_04135_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12118_ (.A1(_04092_),
    .A2(_04132_),
    .B(_04153_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12119_ (.A1(\channels.env_counter[0][13] ),
    .A2(_04135_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12120_ (.A1(_04096_),
    .A2(_04132_),
    .B(_04154_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12121_ (.A1(\channels.env_counter[0][14] ),
    .A2(_04135_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12122_ (.A1(_04100_),
    .A2(_04132_),
    .B(_04155_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12123_ (.A1(_01250_),
    .A2(_03560_),
    .B(_03561_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12124_ (.I0(_03554_),
    .I1(\channels.adsr_state[2][0] ),
    .S(_04156_),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12125_ (.I(_04157_),
    .Z(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12126_ (.I0(_03564_),
    .I1(\channels.adsr_state[2][1] ),
    .S(_04156_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12127_ (.I(_04158_),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12128_ (.A1(_01229_),
    .A2(_03560_),
    .B(_01943_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12129_ (.I0(_03554_),
    .I1(\channels.adsr_state[1][0] ),
    .S(_04159_),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12130_ (.I(_04160_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12131_ (.I0(_03564_),
    .I1(\channels.adsr_state[1][1] ),
    .S(_04159_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12132_ (.I(_04161_),
    .Z(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12133_ (.I(\channels.accum[3][0] ),
    .Z(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12134_ (.I(_04162_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12135_ (.I(\channels.accum[3][1] ),
    .Z(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12136_ (.I(_04163_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12137_ (.I(\channels.accum[3][2] ),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12138_ (.I(_04164_),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12139_ (.I(\channels.accum[3][3] ),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12140_ (.I(_04165_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12141_ (.I(\channels.accum[3][4] ),
    .Z(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12142_ (.I(_04166_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12143_ (.I(\channels.accum[3][5] ),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12144_ (.I(_04167_),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12145_ (.I(\channels.accum[3][6] ),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12146_ (.I(_04168_),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12147_ (.I(\channels.accum[3][7] ),
    .Z(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12148_ (.I(_04169_),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12149_ (.I(\channels.accum[3][8] ),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12150_ (.I(_04170_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12151_ (.I(\channels.accum[3][9] ),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12152_ (.I(_04171_),
    .Z(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12153_ (.I(\channels.accum[3][10] ),
    .Z(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12154_ (.I(_04172_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12155_ (.I(\channels.accum[3][11] ),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12156_ (.I(_04173_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12157_ (.I(\channels.accum[3][12] ),
    .Z(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12158_ (.I(_04174_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12159_ (.I(\channels.accum[3][13] ),
    .Z(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12160_ (.I(_04175_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12161_ (.I(\channels.accum[3][14] ),
    .Z(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12162_ (.I(_04176_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12163_ (.I(\channels.accum[3][15] ),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12164_ (.I(_04177_),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12165_ (.I(\channels.accum[3][16] ),
    .Z(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12166_ (.I(_04178_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12167_ (.I(\channels.accum[3][17] ),
    .Z(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12168_ (.I(_04179_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12169_ (.I(\channels.accum[3][18] ),
    .Z(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12170_ (.I(_04180_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12171_ (.I(\channels.accum[3][19] ),
    .Z(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12172_ (.I(_04181_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12173_ (.I(\channels.accum[3][20] ),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12174_ (.I(_04182_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12175_ (.I(\channels.accum[3][21] ),
    .Z(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12176_ (.I(_04183_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12177_ (.I(\channels.accum[3][22] ),
    .Z(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12178_ (.I(_04184_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12179_ (.I(\channels.accum[3][23] ),
    .Z(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12180_ (.I(_04185_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12181_ (.I(_01104_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12182_ (.A1(_04186_),
    .A2(_03228_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12183_ (.I(_04187_),
    .Z(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12184_ (.I(_04188_),
    .Z(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _12185_ (.A1(_03192_),
    .A2(_03314_),
    .A3(_03198_),
    .A4(\filters.high[5] ),
    .Z(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12186_ (.I(_04190_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12187_ (.I(_04191_),
    .Z(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12188_ (.A1(_03319_),
    .A2(_04192_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _12189_ (.A1(_03182_),
    .A2(_03184_),
    .A3(_03197_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12190_ (.I(net33),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12191_ (.I(_04195_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12192_ (.I(_04196_),
    .Z(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12193_ (.I(_04197_),
    .Z(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12194_ (.A1(\filters.res_lut[3] ),
    .A2(_04198_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12195_ (.A1(_04193_),
    .A2(_04199_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12196_ (.A1(\filters.res_lut[1] ),
    .A2(_04195_),
    .Z(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12197_ (.I(_04201_),
    .Z(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12198_ (.I(_04202_),
    .Z(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12199_ (.I(_04203_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _12200_ (.A1(_03313_),
    .A2(_03314_),
    .A3(_03315_),
    .A4(\filters.high[6] ),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _12201_ (.A1(_03333_),
    .A2(_04205_),
    .Z(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12202_ (.I(_04206_),
    .Z(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12203_ (.I(_04207_),
    .Z(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12204_ (.I(_04208_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12205_ (.I(_04209_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12206_ (.A1(_04204_),
    .A2(_04210_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12207_ (.A1(\filters.res_lut[0] ),
    .A2(_04195_),
    .Z(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _12208_ (.I(_04212_),
    .Z(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12209_ (.I(_04213_),
    .Z(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12210_ (.I(_04214_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12211_ (.I(_03186_),
    .Z(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12212_ (.A1(_03240_),
    .A2(_03205_),
    .A3(_04216_),
    .A4(_03345_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12213_ (.I(_04217_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12214_ (.I(_04218_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12215_ (.A1(_03352_),
    .A2(_04215_),
    .A3(_04219_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _12216_ (.A1(\filters.filter_step[2] ),
    .A2(_03194_),
    .A3(_03197_),
    .A4(\filters.high[3] ),
    .Z(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12217_ (.I(_04221_),
    .Z(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12218_ (.I(net68),
    .Z(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12219_ (.I(_04223_),
    .Z(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _12220_ (.A1(\filters.res_lut[4] ),
    .A2(_04196_),
    .Z(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12221_ (.I(_04225_),
    .Z(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12222_ (.I(_04226_),
    .Z(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12223_ (.I(_04227_),
    .Z(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12224_ (.A1(_03290_),
    .A2(_04224_),
    .A3(_04228_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12225_ (.A1(_04220_),
    .A2(_04229_),
    .Z(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12226_ (.A1(_04220_),
    .A2(_04229_),
    .Z(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12227_ (.A1(_04211_),
    .A2(_04230_),
    .B(_04231_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12228_ (.I(_04210_),
    .Z(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12229_ (.A1(\filters.res_lut[2] ),
    .A2(_04197_),
    .Z(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12230_ (.I(_04234_),
    .Z(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12231_ (.A1(_04233_),
    .A2(_04235_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12232_ (.A1(_04232_),
    .A2(_04236_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12233_ (.I(_04234_),
    .Z(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12234_ (.I(_04238_),
    .Z(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12235_ (.A1(_04233_),
    .A2(_04232_),
    .A3(_04239_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12236_ (.A1(_04200_),
    .A2(_04237_),
    .B(_04240_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12237_ (.I(_04216_),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _12238_ (.I(\filters.high[0] ),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12239_ (.A1(_03241_),
    .A2(_03205_),
    .A3(_04242_),
    .A4(_04243_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12240_ (.I(_04244_),
    .Z(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12241_ (.I(_04194_),
    .Z(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12242_ (.I0(\filters.cutoff_lut[6] ),
    .I1(\filters.res_lut[6] ),
    .S(_04246_),
    .Z(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12243_ (.I(_04247_),
    .Z(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12244_ (.I(_04248_),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12245_ (.I(_04249_),
    .Z(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12246_ (.I(_04250_),
    .Z(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12247_ (.I(_04251_),
    .Z(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12248_ (.A1(_03202_),
    .A2(_04245_),
    .A3(_04252_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _12249_ (.A1(_03313_),
    .A2(_03381_),
    .A3(_03315_),
    .A4(\filters.high[1] ),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12250_ (.I(_04254_),
    .Z(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12251_ (.I(_04255_),
    .Z(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _12252_ (.A1(_04195_),
    .A2(\filters.res_lut[5] ),
    .Z(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12253_ (.I(_04257_),
    .Z(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12254_ (.I(_04258_),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12255_ (.I(_04259_),
    .Z(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12256_ (.I(_04260_),
    .Z(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12257_ (.A1(_03257_),
    .A2(_04256_),
    .A3(_04261_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12258_ (.A1(_04253_),
    .A2(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12259_ (.I(_04248_),
    .Z(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12260_ (.I(_04264_),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12261_ (.I(_04265_),
    .Z(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12262_ (.A1(_03257_),
    .A2(_04256_),
    .A3(_04266_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _12263_ (.I0(\filters.cutoff_lut[7] ),
    .I1(\filters.res_lut[7] ),
    .S(_04246_),
    .Z(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12264_ (.I(net48),
    .Z(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12265_ (.I(_04269_),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _12266_ (.I(_04270_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12267_ (.A1(_03202_),
    .A2(_04245_),
    .A3(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _12268_ (.A1(_03248_),
    .A2(_03285_),
    .A3(_03251_),
    .A4(\filters.high[2] ),
    .Z(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12269_ (.I(_04273_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12270_ (.I(_04274_),
    .Z(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12271_ (.I(_04275_),
    .Z(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12272_ (.A1(_03275_),
    .A2(_04276_),
    .A3(_04261_),
    .Z(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12273_ (.A1(_04267_),
    .A2(_04272_),
    .A3(_04277_),
    .Z(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12274_ (.A1(_04263_),
    .A2(_04278_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12275_ (.A1(_04211_),
    .A2(_04220_),
    .A3(_04229_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12276_ (.A1(_04263_),
    .A2(_04278_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12277_ (.A1(_04279_),
    .A2(_04280_),
    .B(_04281_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12278_ (.A1(_04267_),
    .A2(_04272_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12279_ (.A1(_04267_),
    .A2(_04272_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12280_ (.A1(_04277_),
    .A2(_04283_),
    .B(_04284_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12281_ (.I(_04268_),
    .Z(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12282_ (.I(_04286_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12283_ (.I(_04287_),
    .Z(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12284_ (.A1(_03256_),
    .A2(_04256_),
    .A3(_04288_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12285_ (.A1(_03274_),
    .A2(_04276_),
    .A3(_04265_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12286_ (.A1(_03290_),
    .A2(_04224_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12287_ (.A1(\filters.res_lut[5] ),
    .A2(_04196_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12288_ (.A1(_04291_),
    .A2(_04292_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12289_ (.A1(_04289_),
    .A2(_04290_),
    .A3(_04293_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12290_ (.I(_04202_),
    .Z(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12291_ (.I(_04295_),
    .Z(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12292_ (.A1(_03350_),
    .A2(_04217_),
    .Z(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12293_ (.I(_04297_),
    .Z(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12294_ (.I(_04298_),
    .Z(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12295_ (.A1(_04296_),
    .A2(_04299_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12296_ (.A1(_03241_),
    .A2(_03205_),
    .A3(_04242_),
    .A4(_03361_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12297_ (.A1(_03364_),
    .A2(_04301_),
    .Z(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12298_ (.I(_04302_),
    .Z(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12299_ (.I(_04303_),
    .Z(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12300_ (.I(_04304_),
    .Z(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12301_ (.I(_04213_),
    .Z(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _12302_ (.I(_04306_),
    .Z(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12303_ (.A1(_04305_),
    .A2(_04307_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12304_ (.A1(_03183_),
    .A2(_03184_),
    .A3(_03186_),
    .A4(_03300_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12305_ (.A1(_03303_),
    .A2(_04309_),
    .Z(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12306_ (.I(_04310_),
    .Z(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12307_ (.I(_04311_),
    .Z(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12308_ (.I(_04312_),
    .Z(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12309_ (.A1(_04313_),
    .A2(_04228_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _12310_ (.A1(_04300_),
    .A2(_04308_),
    .A3(_04314_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12311_ (.A1(_04285_),
    .A2(_04294_),
    .A3(_04315_),
    .Z(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12312_ (.A1(_04282_),
    .A2(_04316_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12313_ (.A1(\filters.res_lut[3] ),
    .A2(_04197_),
    .Z(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12314_ (.I(_04318_),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12315_ (.I(_04319_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12316_ (.A1(_04233_),
    .A2(_04320_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12317_ (.I(_04304_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12318_ (.I(_04322_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12319_ (.I(_04215_),
    .Z(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12320_ (.I(_04225_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12321_ (.I(_04325_),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12322_ (.I(_04326_),
    .Z(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12323_ (.A1(_04323_),
    .A2(_04324_),
    .B1(_04327_),
    .B2(_04313_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12324_ (.A1(_04313_),
    .A2(_04322_),
    .A3(_04215_),
    .A4(_04327_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12325_ (.A1(_04300_),
    .A2(_04328_),
    .B(_04329_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12326_ (.I(_04299_),
    .Z(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12327_ (.A1(_04331_),
    .A2(_04238_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12328_ (.A1(_04330_),
    .A2(_04332_),
    .Z(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12329_ (.A1(_04321_),
    .A2(_04333_),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12330_ (.A1(_04317_),
    .A2(_04334_),
    .Z(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12331_ (.A1(_04282_),
    .A2(_04316_),
    .A3(_04334_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12332_ (.A1(_04241_),
    .A2(_04335_),
    .B(_04336_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _12333_ (.I(_04337_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12334_ (.A1(_04241_),
    .A2(_04335_),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12335_ (.A1(_03201_),
    .A2(_04245_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12336_ (.I(_04340_),
    .Z(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12337_ (.I(_04341_),
    .Z(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12338_ (.I0(\filters.cutoff_lut[9] ),
    .I1(\filters.res_lut[9] ),
    .S(net56),
    .Z(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12339_ (.I(_04343_),
    .Z(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12340_ (.I(_04344_),
    .Z(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12341_ (.I(_04345_),
    .Z(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12342_ (.I(_04346_),
    .Z(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12343_ (.A1(_04342_),
    .A2(_04347_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12344_ (.A1(_03255_),
    .A2(_04254_),
    .Z(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12345_ (.I(_04349_),
    .Z(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12346_ (.I(_04350_),
    .Z(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _12347_ (.I0(\filters.cutoff_lut[8] ),
    .I1(\filters.res_lut[8] ),
    .S(net56),
    .Z(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12348_ (.I(_04352_),
    .Z(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12349_ (.I(_04353_),
    .Z(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12350_ (.I(_04354_),
    .Z(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12351_ (.A1(_04351_),
    .A2(_04355_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12352_ (.A1(_04348_),
    .A2(_04356_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12353_ (.A1(_04289_),
    .A2(_04290_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12354_ (.A1(_04289_),
    .A2(_04290_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12355_ (.A1(_04293_),
    .A2(_04358_),
    .B(_04359_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12356_ (.I(_04309_),
    .Z(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12357_ (.A1(_03304_),
    .A2(_04361_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12358_ (.A1(_04292_),
    .A2(_04362_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12359_ (.A1(_03273_),
    .A2(_04286_),
    .A3(_04274_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12360_ (.I(_04247_),
    .Z(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12361_ (.A1(_03289_),
    .A2(_04365_),
    .A3(_04223_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12362_ (.A1(_04364_),
    .A2(_04366_),
    .Z(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12363_ (.A1(_04363_),
    .A2(_04367_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12364_ (.A1(_04360_),
    .A2(_04368_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12365_ (.A1(_04322_),
    .A2(_04296_),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12366_ (.A1(_03240_),
    .A2(_03185_),
    .A3(_04216_),
    .A4(_03375_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12367_ (.I(_04371_),
    .Z(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12368_ (.I(_04212_),
    .Z(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12369_ (.A1(_03385_),
    .A2(_04372_),
    .A3(_04373_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12370_ (.A1(_03318_),
    .A2(_04192_),
    .A3(_04226_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12371_ (.A1(_04374_),
    .A2(_04375_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12372_ (.A1(_04376_),
    .A2(_04370_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12373_ (.I(_04377_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12374_ (.A1(_04369_),
    .A2(_04378_),
    .Z(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12375_ (.A1(_04285_),
    .A2(_04294_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12376_ (.A1(_04285_),
    .A2(_04294_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12377_ (.A1(_04380_),
    .A2(_04315_),
    .B(_04381_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12378_ (.A1(_04357_),
    .A2(_04379_),
    .A3(_04382_),
    .Z(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12379_ (.I(_04342_),
    .Z(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12380_ (.I(_04384_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12381_ (.I(_04355_),
    .Z(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12382_ (.A1(_04385_),
    .A2(_04386_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12383_ (.A1(_04285_),
    .A2(_04294_),
    .A3(_04315_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12384_ (.A1(_04282_),
    .A2(_04388_),
    .Z(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12385_ (.A1(_04387_),
    .A2(_04389_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12386_ (.A1(_04383_),
    .A2(_04390_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12387_ (.A1(_04383_),
    .A2(_04390_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12388_ (.A1(_04339_),
    .A2(_04391_),
    .B(_04392_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12389_ (.A1(_04379_),
    .A2(_04382_),
    .Z(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12390_ (.A1(_04357_),
    .A2(_04394_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12391_ (.A1(_04348_),
    .A2(_04356_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12392_ (.I(_04352_),
    .Z(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12393_ (.I(_04397_),
    .Z(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12394_ (.A1(_03272_),
    .A2(_04274_),
    .Z(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12395_ (.I(_04399_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12396_ (.A1(_04398_),
    .A2(_04400_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12397_ (.A1(_04345_),
    .A2(_04350_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12398_ (.I0(\filters.cutoff_lut[10] ),
    .I1(\filters.res_lut[10] ),
    .S(net34),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12399_ (.I(_04403_),
    .Z(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12400_ (.I(_04404_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12401_ (.I(_04405_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12402_ (.I(_04406_),
    .Z(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12403_ (.A1(_04341_),
    .A2(_04407_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12404_ (.A1(_04401_),
    .A2(_04402_),
    .A3(_04408_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12405_ (.A1(_04396_),
    .A2(_04409_),
    .Z(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12406_ (.A1(_04364_),
    .A2(_04366_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12407_ (.A1(_04363_),
    .A2(_04367_),
    .B(_04411_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _12408_ (.A1(_04190_),
    .A2(_03317_),
    .Z(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12409_ (.I(_04413_),
    .Z(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12410_ (.I(_04414_),
    .Z(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12411_ (.A1(_04415_),
    .A2(_04259_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12412_ (.I(_04286_),
    .Z(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12413_ (.A1(_03288_),
    .A2(_04222_),
    .Z(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12414_ (.I(_04418_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12415_ (.A1(_04417_),
    .A2(_04419_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12416_ (.I(_04264_),
    .Z(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12417_ (.I(_04311_),
    .Z(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12418_ (.A1(_04421_),
    .A2(_04422_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12419_ (.A1(_04416_),
    .A2(_04420_),
    .A3(_04423_),
    .Z(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12420_ (.A1(_03383_),
    .A2(_04371_),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12421_ (.I(_04425_),
    .Z(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12422_ (.I(_04426_),
    .Z(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12423_ (.A1(_04295_),
    .A2(_04427_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12424_ (.A1(_04227_),
    .A2(_04209_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _12425_ (.A1(_03192_),
    .A2(_03314_),
    .A3(_03198_),
    .A4(\filters.high[10] ),
    .Z(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12426_ (.I(_04430_),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12427_ (.A1(_03400_),
    .A2(_04431_),
    .Z(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12428_ (.I(_04432_),
    .Z(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12429_ (.I(_04433_),
    .Z(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12430_ (.A1(_04307_),
    .A2(_04434_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12431_ (.A1(_04428_),
    .A2(_04429_),
    .A3(_04435_),
    .Z(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12432_ (.A1(_04412_),
    .A2(_04424_),
    .A3(_04436_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12433_ (.I(_04437_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12434_ (.A1(_04360_),
    .A2(_04368_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12435_ (.A1(_04369_),
    .A2(_04378_),
    .B(_04439_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12436_ (.A1(_04410_),
    .A2(_04438_),
    .A3(_04440_),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12437_ (.A1(_04369_),
    .A2(net37),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12438_ (.A1(_04442_),
    .A2(_04382_),
    .Z(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12439_ (.A1(_04331_),
    .A2(_04239_),
    .A3(_04330_),
    .Z(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12440_ (.A1(_04321_),
    .A2(_04333_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12441_ (.A1(_04444_),
    .A2(_04445_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12442_ (.I(_04319_),
    .Z(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12443_ (.A1(_04331_),
    .A2(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12444_ (.A1(_04374_),
    .A2(_04375_),
    .Z(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12445_ (.A1(_04370_),
    .A2(_04376_),
    .B(_04449_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12446_ (.A1(_04323_),
    .A2(_04235_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12447_ (.A1(_04450_),
    .A2(_04451_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12448_ (.A1(_04448_),
    .A2(_04452_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12449_ (.A1(_04443_),
    .A2(_04446_),
    .A3(_04453_),
    .Z(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12450_ (.A1(_04395_),
    .A2(_04441_),
    .A3(_04454_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12451_ (.A1(_04393_),
    .A2(_04455_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12452_ (.A1(_04393_),
    .A2(_04455_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _12453_ (.A1(_04338_),
    .A2(_04456_),
    .B(_04457_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12454_ (.I(_04443_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12455_ (.A1(_04443_),
    .A2(_04453_),
    .Z(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12456_ (.A1(_04446_),
    .A2(_04460_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12457_ (.A1(_04459_),
    .A2(_04453_),
    .B(_04461_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12458_ (.A1(_04357_),
    .A2(_04394_),
    .B(_04441_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _12459_ (.A1(_04357_),
    .A2(_04394_),
    .A3(_04441_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12460_ (.A1(_04463_),
    .A2(_04454_),
    .B(_04464_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12461_ (.A1(_04437_),
    .A2(_04440_),
    .Z(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12462_ (.A1(_04410_),
    .A2(_04466_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _12463_ (.A1(\filters.filter_step[2] ),
    .A2(_03184_),
    .A3(\filters.filter_step[0] ),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12464_ (.I(_04468_),
    .Z(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12465_ (.A1(\filters.cutoff_lut[11] ),
    .A2(_04469_),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12466_ (.I(_04470_),
    .Z(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12467_ (.I(_04471_),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12468_ (.I(_04472_),
    .Z(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12469_ (.I(_04473_),
    .Z(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12470_ (.I(_04474_),
    .Z(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12471_ (.A1(_04384_),
    .A2(_04475_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12472_ (.I(_04345_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12473_ (.I(_04404_),
    .Z(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12474_ (.I(_04478_),
    .Z(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12475_ (.I(_04479_),
    .Z(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12476_ (.I(_04480_),
    .Z(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12477_ (.A1(_04477_),
    .A2(_04351_),
    .B1(_04481_),
    .B2(_04341_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12478_ (.A1(_04341_),
    .A2(_04477_),
    .A3(_04350_),
    .A4(_04407_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12479_ (.A1(_04401_),
    .A2(_04482_),
    .B(_04483_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12480_ (.A1(_04397_),
    .A2(_04419_),
    .Z(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12481_ (.A1(_03256_),
    .A2(_04255_),
    .A3(_04405_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12482_ (.A1(_03275_),
    .A2(_04345_),
    .A3(_04276_),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12483_ (.A1(_04485_),
    .A2(_04486_),
    .A3(_04487_),
    .Z(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12484_ (.A1(_04484_),
    .A2(_04488_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12485_ (.A1(_04476_),
    .A2(_04489_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12486_ (.A1(_04412_),
    .A2(_04424_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12487_ (.A1(_04412_),
    .A2(_04424_),
    .Z(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12488_ (.A1(_04491_),
    .A2(_04436_),
    .B(_04492_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _12489_ (.A1(_04348_),
    .A2(_04356_),
    .A3(_04409_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12490_ (.I(_04287_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12491_ (.I(_04419_),
    .Z(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12492_ (.I(_04311_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _12493_ (.A1(_04495_),
    .A2(_04496_),
    .B1(_04497_),
    .B2(_04250_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12494_ (.A1(_04495_),
    .A2(_04250_),
    .A3(_04419_),
    .A4(_04497_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12495_ (.A1(net60),
    .A2(_04498_),
    .B(_04499_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12496_ (.I(_04257_),
    .Z(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12497_ (.I(_04206_),
    .Z(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12498_ (.A1(_04501_),
    .A2(_04502_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12499_ (.I(_04310_),
    .Z(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12500_ (.A1(_04269_),
    .A2(_04504_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12501_ (.I(_04365_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12502_ (.I(_04414_),
    .Z(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12503_ (.A1(_04506_),
    .A2(_04507_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _12504_ (.A1(_04503_),
    .A2(_04505_),
    .A3(_04508_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12505_ (.A1(_04202_),
    .A2(_04433_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12506_ (.I(_04297_),
    .Z(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12507_ (.A1(_04226_),
    .A2(_04511_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12508_ (.I(_04373_),
    .Z(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12509_ (.A1(_03240_),
    .A2(_03185_),
    .A3(_04216_),
    .A4(_03412_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12510_ (.A1(_03415_),
    .A2(_04514_),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12511_ (.I(_04515_),
    .Z(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12512_ (.I(_04516_),
    .Z(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12513_ (.A1(_04513_),
    .A2(_04517_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12514_ (.A1(_04510_),
    .A2(_04512_),
    .A3(_04518_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12515_ (.A1(_04500_),
    .A2(_04509_),
    .A3(net67),
    .Z(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12516_ (.A1(_04494_),
    .A2(_04520_),
    .Z(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12517_ (.A1(_04490_),
    .A2(_04493_),
    .A3(_04521_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12518_ (.A1(_04438_),
    .A2(_04440_),
    .Z(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12519_ (.I(_04239_),
    .Z(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12520_ (.A1(_04323_),
    .A2(_04524_),
    .A3(_04450_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12521_ (.I(_04320_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12522_ (.A1(_04331_),
    .A2(_04526_),
    .A3(_04452_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12523_ (.A1(_04525_),
    .A2(_04527_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12524_ (.A1(_04323_),
    .A2(_04320_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12525_ (.I(_04228_),
    .Z(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12526_ (.I(_04434_),
    .Z(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12527_ (.I(_04531_),
    .Z(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12528_ (.A1(_04530_),
    .A2(_04233_),
    .B1(_04532_),
    .B2(_04324_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _12529_ (.A1(_04324_),
    .A2(_04327_),
    .A3(_04210_),
    .A4(_04532_),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12530_ (.A1(_04428_),
    .A2(_04533_),
    .B(_04534_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12531_ (.I(_04426_),
    .Z(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12532_ (.I(_04536_),
    .Z(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12533_ (.I(_04537_),
    .Z(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12534_ (.A1(_04538_),
    .A2(_04238_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12535_ (.A1(_04535_),
    .A2(_04539_),
    .Z(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12536_ (.A1(_04529_),
    .A2(_04540_),
    .Z(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12537_ (.A1(_04523_),
    .A2(_04528_),
    .A3(_04541_),
    .Z(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12538_ (.A1(_04467_),
    .A2(_04522_),
    .A3(_04542_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12539_ (.A1(_04543_),
    .A2(_04465_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12540_ (.A1(_04462_),
    .A2(_04544_),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12541_ (.A1(_04458_),
    .A2(_04545_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12542_ (.A1(_04253_),
    .A2(_04262_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12543_ (.I(_04205_),
    .Z(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12544_ (.A1(_03335_),
    .A2(_04324_),
    .A3(_04548_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12545_ (.A1(_03275_),
    .A2(_04276_),
    .A3(_04327_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12546_ (.I(_04296_),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12547_ (.A1(_03319_),
    .A2(_04551_),
    .A3(_04192_),
    .Z(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12548_ (.A1(_04549_),
    .A2(_04550_),
    .A3(_04552_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12549_ (.A1(_04547_),
    .A2(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12550_ (.I(_04203_),
    .Z(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12551_ (.A1(_03335_),
    .A2(_04555_),
    .A3(_04548_),
    .Z(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12552_ (.A1(_04556_),
    .A2(_04220_),
    .A3(_04229_),
    .Z(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12553_ (.A1(_04263_),
    .A2(_04278_),
    .A3(_04557_),
    .Z(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12554_ (.A1(_04558_),
    .A2(_04554_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12555_ (.A1(_04200_),
    .A2(_04237_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12556_ (.A1(_04362_),
    .A2(_04199_),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12557_ (.A1(\filters.res_lut[1] ),
    .A2(_04196_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12558_ (.A1(_04549_),
    .A2(_04550_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12559_ (.A1(_04549_),
    .A2(_04550_),
    .Z(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _12560_ (.A1(_04562_),
    .A2(_04193_),
    .A3(_04563_),
    .B(_04564_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12561_ (.A1(\filters.res_lut[2] ),
    .A2(_04197_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12562_ (.A1(_04193_),
    .A2(_04566_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12563_ (.A1(_04565_),
    .A2(_04567_),
    .Z(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12564_ (.A1(_04565_),
    .A2(_04567_),
    .Z(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12565_ (.A1(_04561_),
    .A2(_04568_),
    .B(_04569_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12566_ (.A1(_04200_),
    .A2(_04237_),
    .A3(_04559_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _12567_ (.A1(_04570_),
    .A2(_04571_),
    .Z(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12568_ (.A1(_04559_),
    .A2(_04560_),
    .B(_04572_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12569_ (.A1(_04387_),
    .A2(_04282_),
    .A3(net47),
    .Z(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12570_ (.A1(_04570_),
    .A2(_04571_),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12571_ (.A1(_04574_),
    .A2(_04572_),
    .A3(_04575_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12572_ (.A1(_04317_),
    .A2(_04241_),
    .A3(_04334_),
    .Z(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12573_ (.A1(_04383_),
    .A2(_04390_),
    .A3(_04577_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12574_ (.A1(_04576_),
    .A2(_04578_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12575_ (.A1(_04576_),
    .A2(_04578_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12576_ (.A1(_04573_),
    .A2(_04579_),
    .B(_04580_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12577_ (.A1(_04393_),
    .A2(_04455_),
    .A3(_04338_),
    .Z(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12578_ (.A1(_04581_),
    .A2(_04582_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12579_ (.A1(_04574_),
    .A2(_04570_),
    .A3(_04571_),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12580_ (.A1(_04554_),
    .A2(_04558_),
    .Z(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12581_ (.I(_04447_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12582_ (.I(_04586_),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12583_ (.A1(_04496_),
    .A2(_04587_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12584_ (.A1(_04362_),
    .A2(_04562_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12585_ (.I(_04215_),
    .Z(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12586_ (.A1(_03319_),
    .A2(_04590_),
    .A3(_04192_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12587_ (.I(_04256_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12588_ (.A1(_03257_),
    .A2(_04592_),
    .A3(_04530_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12589_ (.A1(_04591_),
    .A2(_04593_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12590_ (.A1(_04591_),
    .A2(_04593_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12591_ (.A1(_04589_),
    .A2(_04594_),
    .B(_04595_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12592_ (.I(_04313_),
    .Z(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12593_ (.A1(_04597_),
    .A2(_04524_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12594_ (.A1(_04596_),
    .A2(_04598_),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12595_ (.A1(_04596_),
    .A2(_04598_),
    .Z(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12596_ (.A1(_04588_),
    .A2(_04599_),
    .B(_04600_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12597_ (.I(_04261_),
    .Z(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12598_ (.I(_04602_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12599_ (.I(_04603_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12600_ (.A1(_04385_),
    .A2(_04604_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12601_ (.I(_04551_),
    .Z(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12602_ (.A1(_03304_),
    .A2(_04361_),
    .A3(_04606_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12603_ (.A1(_04591_),
    .A2(_04593_),
    .A3(_04607_),
    .Z(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12604_ (.A1(_04605_),
    .A2(_04608_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12605_ (.A1(_04547_),
    .A2(_04553_),
    .Z(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12606_ (.A1(_04609_),
    .A2(_04610_),
    .Z(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12607_ (.A1(_04565_),
    .A2(_04567_),
    .A3(_04561_),
    .Z(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12608_ (.A1(_04611_),
    .A2(_04612_),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12609_ (.A1(_04601_),
    .A2(_04613_),
    .Z(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12610_ (.A1(_04584_),
    .A2(_04585_),
    .A3(_04614_),
    .Z(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12611_ (.A1(_04601_),
    .A2(_04613_),
    .Z(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12612_ (.A1(_04611_),
    .A2(_04612_),
    .B(_04616_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12613_ (.A1(_04585_),
    .A2(_04614_),
    .B(_04584_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _12614_ (.A1(_04615_),
    .A2(_04617_),
    .A3(_04618_),
    .Z(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12615_ (.A1(_04609_),
    .A2(_04610_),
    .Z(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12616_ (.A1(_03274_),
    .A2(_04275_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12617_ (.I(_04621_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12618_ (.A1(_04622_),
    .A2(_04199_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12619_ (.I(_04555_),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12620_ (.I(_04624_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12621_ (.A1(_04496_),
    .A2(_04625_),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12622_ (.I(_04590_),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12623_ (.I(_04530_),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12624_ (.I(_04628_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12625_ (.A1(_04597_),
    .A2(_04627_),
    .B1(_04629_),
    .B2(_04384_),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12626_ (.A1(_04384_),
    .A2(_04597_),
    .A3(_04627_),
    .A4(_04628_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12627_ (.A1(_04626_),
    .A2(_04630_),
    .B(_04631_),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12628_ (.A1(_04291_),
    .A2(_04566_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12629_ (.A1(_04632_),
    .A2(_04633_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12630_ (.A1(_04632_),
    .A2(_04633_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12631_ (.A1(_04623_),
    .A2(_04634_),
    .B(_04635_),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12632_ (.A1(_04588_),
    .A2(_04599_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12633_ (.A1(_04620_),
    .A2(_04636_),
    .A3(_04637_),
    .Z(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12634_ (.A1(_04605_),
    .A2(_04608_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12635_ (.I(_04639_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12636_ (.A1(_03258_),
    .A2(_04592_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12637_ (.A1(_04641_),
    .A2(_04199_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12638_ (.I(_04400_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12639_ (.I(_04606_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12640_ (.I(_04644_),
    .Z(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12641_ (.I(_04590_),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12642_ (.A1(_04643_),
    .A2(_04496_),
    .A3(_04645_),
    .A4(_04646_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12643_ (.I(_04524_),
    .Z(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12644_ (.A1(_04643_),
    .A2(_04648_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12645_ (.A1(_04647_),
    .A2(_04649_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12646_ (.A1(_04566_),
    .A2(_04647_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12647_ (.A1(_04642_),
    .A2(_04650_),
    .B(_04651_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12648_ (.A1(_04632_),
    .A2(_04633_),
    .A3(_04623_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12649_ (.A1(_04652_),
    .A2(_04653_),
    .Z(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12650_ (.A1(_04652_),
    .A2(_04653_),
    .Z(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12651_ (.A1(_04640_),
    .A2(_04654_),
    .B(_04655_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12652_ (.I(_04385_),
    .Z(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12653_ (.I(_04447_),
    .Z(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12654_ (.I(_04658_),
    .Z(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12655_ (.I(_04659_),
    .Z(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12656_ (.I(_04648_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12657_ (.I(_04645_),
    .Z(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _12658_ (.A1(_03258_),
    .A2(_04592_),
    .A3(_04662_),
    .A4(_04646_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12659_ (.A1(_04643_),
    .A2(_04661_),
    .A3(_04663_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12660_ (.I(_04646_),
    .Z(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12661_ (.A1(_03258_),
    .A2(_04592_),
    .A3(_04662_),
    .A4(_04665_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _12662_ (.A1(_04641_),
    .A2(_04566_),
    .B1(_04666_),
    .B2(_04622_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _12663_ (.A1(_04657_),
    .A2(_04660_),
    .A3(_04664_),
    .A4(_04667_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12664_ (.I(_04587_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _12665_ (.A1(_04657_),
    .A2(_04669_),
    .B1(_04664_),
    .B2(_04667_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12666_ (.I(_04234_),
    .Z(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12667_ (.I(_04671_),
    .Z(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12668_ (.I(_04672_),
    .Z(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _12669_ (.I(_04673_),
    .Z(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12670_ (.I(_04674_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _12671_ (.A1(_04657_),
    .A2(_04675_),
    .A3(_04663_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12672_ (.A1(_04668_),
    .A2(_04670_),
    .B(_04676_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12673_ (.A1(\filters.res_lut[0] ),
    .A2(_04198_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _12674_ (.A1(_04622_),
    .A2(_04562_),
    .B1(_04678_),
    .B2(_04291_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12675_ (.A1(_04647_),
    .A2(_04679_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _12676_ (.A1(_04668_),
    .A2(_04670_),
    .A3(_04676_),
    .B(_04680_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12677_ (.A1(_04677_),
    .A2(_04681_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12678_ (.A1(_04597_),
    .A2(_04665_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12679_ (.A1(_04385_),
    .A2(_04629_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _12680_ (.A1(_04683_),
    .A2(_04684_),
    .A3(_04626_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12681_ (.I0(_04674_),
    .I1(_04649_),
    .S(_04647_),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12682_ (.A1(_04642_),
    .A2(_04686_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12683_ (.I(_04664_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _12684_ (.A1(_04688_),
    .A2(_04668_),
    .Z(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12685_ (.A1(_04685_),
    .A2(_04687_),
    .A3(_04689_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12686_ (.A1(_04652_),
    .A2(_04653_),
    .A3(_04640_),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12687_ (.A1(_04682_),
    .A2(_04690_),
    .B(_04691_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _12688_ (.A1(_04685_),
    .A2(_04687_),
    .A3(_04689_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _12689_ (.A1(_04668_),
    .A2(_04670_),
    .B(_04676_),
    .C(_04680_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12690_ (.A1(_04351_),
    .A2(_04662_),
    .B1(_04665_),
    .B2(_04643_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12691_ (.A1(_04622_),
    .A2(_04666_),
    .B(_04657_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12692_ (.I(_04661_),
    .Z(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12693_ (.A1(_04697_),
    .A2(_04663_),
    .B(_04676_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _12694_ (.A1(_04695_),
    .A2(_04696_),
    .A3(_04698_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _12695_ (.A1(_04677_),
    .A2(_04681_),
    .B1(_04694_),
    .B2(_04699_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12696_ (.A1(_04687_),
    .A2(_04689_),
    .B(_04685_),
    .ZN(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12697_ (.A1(_04687_),
    .A2(_04689_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _12698_ (.A1(_04693_),
    .A2(_04700_),
    .B(_04701_),
    .C(_04702_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _12699_ (.A1(_04638_),
    .A2(_04656_),
    .B1(_04692_),
    .B2(_04703_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12700_ (.A1(_04638_),
    .A2(_04656_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12701_ (.I(_04585_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12702_ (.A1(_04706_),
    .A2(_04614_),
    .Z(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12703_ (.A1(_04704_),
    .A2(_04705_),
    .B(_04707_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12704_ (.A1(_04636_),
    .A2(_04637_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12705_ (.A1(_04636_),
    .A2(_04637_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12706_ (.A1(_04620_),
    .A2(_04709_),
    .B(_04710_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _12707_ (.A1(_04707_),
    .A2(_04704_),
    .A3(_04705_),
    .B(_04711_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12708_ (.A1(_04615_),
    .A2(_04618_),
    .B(_04617_),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12709_ (.A1(_04619_),
    .A2(_04708_),
    .A3(_04712_),
    .A4(_04713_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12710_ (.A1(_04576_),
    .A2(_04578_),
    .A3(_04573_),
    .Z(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12711_ (.A1(_04584_),
    .A2(_04585_),
    .A3(_04614_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12712_ (.A1(_04617_),
    .A2(_04618_),
    .B(_04716_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12713_ (.A1(_04715_),
    .A2(_04717_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12714_ (.A1(_04715_),
    .A2(_04717_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12715_ (.A1(_04714_),
    .A2(_04718_),
    .B(_04719_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12716_ (.A1(_04581_),
    .A2(_04582_),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _12717_ (.A1(_04458_),
    .A2(_04545_),
    .B1(_04583_),
    .B2(_04720_),
    .C(_04721_),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _12718_ (.A1(_04546_),
    .A2(_04722_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12719_ (.I(_04495_),
    .Z(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12720_ (.I(_04414_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12721_ (.I(_04725_),
    .Z(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _12722_ (.A1(_04724_),
    .A2(_04312_),
    .B1(_04726_),
    .B2(_04251_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12723_ (.I(_04288_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _12724_ (.A1(_04728_),
    .A2(_04251_),
    .A3(_04312_),
    .A4(_04726_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _12725_ (.A1(_04503_),
    .A2(_04727_),
    .B(_04729_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12726_ (.A1(_04417_),
    .A2(_04507_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12727_ (.I(_04248_),
    .Z(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12728_ (.A1(_04732_),
    .A2(_04208_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12729_ (.I(_04501_),
    .Z(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12730_ (.A1(_04734_),
    .A2(_04298_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12731_ (.A1(_04731_),
    .A2(_04733_),
    .A3(_04735_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12732_ (.A1(_04730_),
    .A2(_04736_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12733_ (.A1(_04295_),
    .A2(_04517_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12734_ (.I(_03187_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12735_ (.I0(\filters.high[12] ),
    .I1(\filters.band[12] ),
    .S(_04739_),
    .Z(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12736_ (.I(_04740_),
    .Z(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12737_ (.I(_04741_),
    .Z(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12738_ (.A1(_04214_),
    .A2(_04742_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12739_ (.A1(_04305_),
    .A2(_04326_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12740_ (.A1(_04738_),
    .A2(_04743_),
    .A3(_04744_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12741_ (.I(_04745_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12742_ (.A1(_04730_),
    .A2(_04736_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12743_ (.A1(_04737_),
    .A2(_04746_),
    .B(_04747_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12744_ (.A1(_04397_),
    .A2(_04504_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12745_ (.A1(_03273_),
    .A2(_04274_),
    .A3(_04405_),
    .Z(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12746_ (.I(_04343_),
    .Z(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12747_ (.I(_04751_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _12748_ (.A1(_03290_),
    .A2(_04752_),
    .A3(_04224_),
    .Z(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12749_ (.A1(_04749_),
    .A2(_04750_),
    .A3(_04753_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12750_ (.A1(_04486_),
    .A2(_04487_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12751_ (.A1(_04486_),
    .A2(_04487_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12752_ (.A1(_04485_),
    .A2(_04755_),
    .B(_04756_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12753_ (.A1(_04754_),
    .A2(_04757_),
    .ZN(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12754_ (.I(_04269_),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12755_ (.I(_04502_),
    .Z(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12756_ (.A1(_04759_),
    .A2(_04725_),
    .B1(_04760_),
    .B2(_04265_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12757_ (.A1(_04759_),
    .A2(_04265_),
    .A3(_04725_),
    .A4(_04760_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12758_ (.A1(_04735_),
    .A2(_04761_),
    .B(_04762_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12759_ (.A1(_04258_),
    .A2(_04302_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12760_ (.A1(_04286_),
    .A2(_04207_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12761_ (.A1(_04264_),
    .A2(_04511_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12762_ (.A1(_04764_),
    .A2(_04765_),
    .A3(_04766_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12763_ (.I(_04740_),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12764_ (.A1(_04201_),
    .A2(_04768_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12765_ (.I0(\filters.high[13] ),
    .I1(\filters.band[13] ),
    .S(_04739_),
    .Z(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12766_ (.I(_04770_),
    .Z(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12767_ (.A1(_04213_),
    .A2(_04771_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12768_ (.A1(_04536_),
    .A2(_04325_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12769_ (.A1(_04769_),
    .A2(_04772_),
    .A3(_04773_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12770_ (.A1(_04763_),
    .A2(_04767_),
    .A3(_04774_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12771_ (.A1(_04775_),
    .A2(_04758_),
    .Z(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12772_ (.A1(_04758_),
    .A2(_04775_),
    .Z(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12773_ (.A1(_04748_),
    .A2(_04776_),
    .B(_04777_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12774_ (.I(_04778_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12775_ (.I(_04515_),
    .Z(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12776_ (.I(_04780_),
    .Z(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12777_ (.I(_04781_),
    .Z(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12778_ (.I(_04782_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12779_ (.A1(_04318_),
    .A2(_04783_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12780_ (.A1(_04772_),
    .A2(_04773_),
    .Z(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12781_ (.A1(_04772_),
    .A2(_04773_),
    .Z(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12782_ (.A1(_04769_),
    .A2(_04785_),
    .B(_04786_),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12783_ (.I(_04742_),
    .Z(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12784_ (.I(_04788_),
    .Z(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12785_ (.A1(_04671_),
    .A2(_04789_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12786_ (.A1(_04784_),
    .A2(_04787_),
    .A3(_04790_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12787_ (.A1(_04779_),
    .A2(_04791_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12788_ (.I(_04532_),
    .Z(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12789_ (.A1(_04319_),
    .A2(_04793_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12790_ (.I(_04235_),
    .Z(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12791_ (.I(_04795_),
    .Z(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12792_ (.I(_04796_),
    .Z(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12793_ (.I(_04517_),
    .Z(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12794_ (.I(_04798_),
    .Z(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12795_ (.A1(_04743_),
    .A2(_04744_),
    .Z(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12796_ (.A1(_04743_),
    .A2(_04744_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12797_ (.A1(_04738_),
    .A2(_04800_),
    .B(_04801_),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12798_ (.A1(_04797_),
    .A2(_04799_),
    .B(_04802_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12799_ (.A1(_04797_),
    .A2(_04799_),
    .A3(_04802_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12800_ (.A1(_04794_),
    .A2(_04803_),
    .B(_04804_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12801_ (.A1(_04778_),
    .A2(_04791_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12802_ (.A1(_04805_),
    .A2(_04806_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12803_ (.A1(_04792_),
    .A2(_04807_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12804_ (.I(_04469_),
    .Z(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12805_ (.A1(\filters.cutoff_lut[11] ),
    .A2(_04809_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12806_ (.A1(_04621_),
    .A2(_04810_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12807_ (.A1(\filters.cutoff_lut[13] ),
    .A2(_04469_),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12808_ (.I(_04812_),
    .Z(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12809_ (.I(_04813_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12810_ (.A1(_03202_),
    .A2(_04245_),
    .A3(_04814_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12811_ (.A1(\filters.cutoff_lut[12] ),
    .A2(_04469_),
    .Z(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12812_ (.I(_04816_),
    .Z(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12813_ (.A1(_03255_),
    .A2(_04255_),
    .A3(_04817_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12814_ (.A1(_04815_),
    .A2(_04818_),
    .Z(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12815_ (.A1(_04811_),
    .A2(_04819_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12816_ (.A1(_04750_),
    .A2(_04753_),
    .Z(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12817_ (.A1(_04750_),
    .A2(_04753_),
    .Z(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12818_ (.A1(_04749_),
    .A2(_04821_),
    .B(_04822_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12819_ (.I(_04470_),
    .Z(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12820_ (.I(_04816_),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _12821_ (.A1(_04340_),
    .A2(_04350_),
    .A3(_04824_),
    .A4(_04825_),
    .Z(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12822_ (.A1(_03317_),
    .A2(_04352_),
    .A3(net58),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12823_ (.A1(net69),
    .A2(net68),
    .A3(_04403_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12824_ (.A1(_03303_),
    .A2(_04343_),
    .A3(_04309_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _12825_ (.A1(_04827_),
    .A2(_04828_),
    .A3(_04829_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12826_ (.A1(_04826_),
    .A2(_04830_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12827_ (.A1(_04823_),
    .A2(_04831_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12828_ (.A1(_04832_),
    .A2(_04820_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12829_ (.I(_04816_),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12830_ (.I(_04834_),
    .Z(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12831_ (.I(_04835_),
    .Z(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12832_ (.I(_04836_),
    .Z(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _12833_ (.A1(_04351_),
    .A2(_04473_),
    .B1(_04837_),
    .B2(_04342_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12834_ (.A1(_04826_),
    .A2(_04838_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12835_ (.A1(_04754_),
    .A2(_04757_),
    .Z(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12836_ (.A1(_04839_),
    .A2(_04840_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12837_ (.A1(_04841_),
    .A2(_04833_),
    .Z(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12838_ (.A1(_04748_),
    .A2(_04776_),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12839_ (.A1(_04833_),
    .A2(_04839_),
    .A3(_04840_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12840_ (.A1(_04842_),
    .A2(net66),
    .B(_04844_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12841_ (.A1(_04820_),
    .A2(_04832_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12842_ (.A1(\filters.cutoff_lut[14] ),
    .A2(_04468_),
    .Z(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12843_ (.I(_04847_),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12844_ (.I(_04848_),
    .Z(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12845_ (.I(_04849_),
    .Z(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12846_ (.I(_04850_),
    .Z(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12847_ (.A1(_04342_),
    .A2(_04851_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12848_ (.A1(_03289_),
    .A2(_04224_),
    .A3(_04824_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12849_ (.A1(_03273_),
    .A2(_04275_),
    .A3(_04817_),
    .ZN(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12850_ (.I(_04813_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12851_ (.I(_04855_),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12852_ (.A1(_03256_),
    .A2(_04255_),
    .A3(_04856_),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12853_ (.A1(_04853_),
    .A2(_04854_),
    .A3(_04857_),
    .Z(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12854_ (.A1(_04852_),
    .A2(_04858_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12855_ (.A1(_04828_),
    .A2(_04829_),
    .Z(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12856_ (.A1(_04828_),
    .A2(_04829_),
    .Z(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _12857_ (.A1(_04827_),
    .A2(_04860_),
    .B(_04861_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12858_ (.A1(_04815_),
    .A2(_04818_),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12859_ (.A1(_04811_),
    .A2(_04819_),
    .B(_04863_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12860_ (.A1(_04353_),
    .A2(_04760_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12861_ (.A1(_04752_),
    .A2(_04507_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12862_ (.A1(_04422_),
    .A2(_04406_),
    .ZN(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12863_ (.A1(_04865_),
    .A2(_04866_),
    .A3(_04867_),
    .Z(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12864_ (.A1(_04862_),
    .A2(_04864_),
    .A3(_04868_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12865_ (.A1(_04859_),
    .A2(_04869_),
    .Z(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12866_ (.A1(_04846_),
    .A2(_04870_),
    .Z(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12867_ (.A1(_04763_),
    .A2(_04767_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12868_ (.I(_04774_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12869_ (.A1(_04763_),
    .A2(_04767_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12870_ (.A1(_04872_),
    .A2(_04873_),
    .B(_04874_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12871_ (.A1(_04826_),
    .A2(_04830_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12872_ (.A1(_04823_),
    .A2(_04831_),
    .B(_04876_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12873_ (.I(_04506_),
    .Z(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12874_ (.I(_04270_),
    .Z(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _12875_ (.A1(_04878_),
    .A2(_04299_),
    .B1(_04209_),
    .B2(_04879_),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12876_ (.I(_04732_),
    .Z(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12877_ (.A1(_04879_),
    .A2(_04881_),
    .A3(_04298_),
    .A4(_04209_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12878_ (.A1(_04764_),
    .A2(_04880_),
    .B(_04882_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12879_ (.A1(_04501_),
    .A2(_04426_),
    .Z(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12880_ (.I(_04301_),
    .Z(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12881_ (.A1(_03365_),
    .A2(_04365_),
    .A3(_04885_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12882_ (.A1(_03351_),
    .A2(_04417_),
    .A3(_04219_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12883_ (.A1(_04884_),
    .A2(_04886_),
    .A3(_04887_),
    .Z(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12884_ (.I(_04770_),
    .Z(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12885_ (.A1(_04202_),
    .A2(_04889_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12886_ (.I0(\filters.high[14] ),
    .I1(\filters.band[14] ),
    .S(_04739_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12887_ (.I(_04891_),
    .Z(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12888_ (.I(_04892_),
    .Z(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12889_ (.A1(_04373_),
    .A2(_04893_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12890_ (.A1(_04227_),
    .A2(_04434_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12891_ (.A1(_04890_),
    .A2(_04894_),
    .A3(_04895_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12892_ (.A1(_04883_),
    .A2(_04888_),
    .A3(_04896_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12893_ (.A1(_04877_),
    .A2(_04897_),
    .Z(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12894_ (.A1(_04875_),
    .A2(_04898_),
    .Z(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12895_ (.A1(_04871_),
    .A2(_04899_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12896_ (.A1(_04845_),
    .A2(_04900_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12897_ (.A1(_04805_),
    .A2(_04806_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12898_ (.A1(_04845_),
    .A2(_04900_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12899_ (.A1(_04901_),
    .A2(_04902_),
    .B(_04903_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12900_ (.A1(_04846_),
    .A2(_04870_),
    .Z(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12901_ (.A1(_04871_),
    .A2(_04899_),
    .B(_04905_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12902_ (.A1(_04859_),
    .A2(_04869_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12903_ (.A1(_04852_),
    .A2(_04858_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _12904_ (.A1(\filters.cutoff_lut[15] ),
    .A2(_04468_),
    .Z(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _12905_ (.I(_04909_),
    .Z(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12906_ (.I(_04910_),
    .Z(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12907_ (.I(_04911_),
    .Z(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12908_ (.A1(_03201_),
    .A2(_04244_),
    .A3(_04912_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12909_ (.I(_04847_),
    .Z(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12910_ (.A1(_03255_),
    .A2(_04254_),
    .A3(_04914_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _12911_ (.A1(_04913_),
    .A2(_04915_),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12912_ (.A1(_03304_),
    .A2(_04361_),
    .A3(_04471_),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12913_ (.A1(_03289_),
    .A2(_04223_),
    .A3(_04834_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12914_ (.A1(_03274_),
    .A2(_04275_),
    .A3(_04855_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12915_ (.A1(_04917_),
    .A2(_04918_),
    .A3(_04919_),
    .Z(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12916_ (.A1(_04916_),
    .A2(_04920_),
    .Z(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _12917_ (.A1(_04346_),
    .A2(_04726_),
    .B1(_04407_),
    .B2(_04312_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _12918_ (.A1(_04346_),
    .A2(_04497_),
    .A3(_04726_),
    .A4(_04480_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _12919_ (.A1(_04865_),
    .A2(_04922_),
    .B(_04923_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12920_ (.I(_04810_),
    .Z(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12921_ (.A1(_04291_),
    .A2(_04925_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12922_ (.A1(_04854_),
    .A2(_04857_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12923_ (.A1(_04854_),
    .A2(_04857_),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _12924_ (.A1(_04926_),
    .A2(_04927_),
    .B(_04928_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12925_ (.A1(_04398_),
    .A2(_04298_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12926_ (.A1(_03334_),
    .A2(_04344_),
    .A3(net70),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _12927_ (.A1(_03318_),
    .A2(_04191_),
    .A3(_04478_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12928_ (.A1(_04931_),
    .A2(_04932_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12929_ (.A1(_04930_),
    .A2(_04933_),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12930_ (.A1(_04924_),
    .A2(_04929_),
    .A3(_04934_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12931_ (.A1(_04908_),
    .A2(_04921_),
    .A3(_04935_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12932_ (.A1(_04883_),
    .A2(_04888_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12933_ (.I(_04896_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12934_ (.A1(_04883_),
    .A2(_04888_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12935_ (.A1(_04937_),
    .A2(_04938_),
    .B(_04939_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12936_ (.A1(_04864_),
    .A2(_04868_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12937_ (.A1(_04864_),
    .A2(_04868_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12938_ (.A1(_04862_),
    .A2(_04941_),
    .B(_04942_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12939_ (.A1(_04886_),
    .A2(_04887_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12940_ (.A1(_04886_),
    .A2(_04887_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12941_ (.A1(_04884_),
    .A2(_04944_),
    .B(_04945_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12942_ (.A1(_04259_),
    .A2(_04433_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12943_ (.A1(_04249_),
    .A2(_04536_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12944_ (.A1(_04759_),
    .A2(_04303_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12945_ (.A1(_04947_),
    .A2(_04948_),
    .A3(_04949_),
    .Z(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12946_ (.A1(_04946_),
    .A2(_04950_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12947_ (.I(_04893_),
    .Z(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12948_ (.A1(_04203_),
    .A2(_04952_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12949_ (.I0(\filters.high[15] ),
    .I1(\filters.band[15] ),
    .S(_03188_),
    .Z(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12950_ (.I(_04954_),
    .Z(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12951_ (.A1(_04513_),
    .A2(_04955_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12952_ (.A1(_04326_),
    .A2(_04798_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _12953_ (.A1(_04953_),
    .A2(_04956_),
    .A3(_04957_),
    .Z(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12954_ (.A1(_04951_),
    .A2(_04958_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _12955_ (.A1(_04940_),
    .A2(_04943_),
    .A3(_04959_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12956_ (.A1(_04907_),
    .A2(_04936_),
    .A3(_04960_),
    .Z(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12957_ (.A1(_04906_),
    .A2(_04961_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12958_ (.A1(_04661_),
    .A2(_04789_),
    .B(_04787_),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12959_ (.A1(_04674_),
    .A2(_04789_),
    .A3(_04787_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12960_ (.A1(_04784_),
    .A2(_04963_),
    .B(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12961_ (.A1(_04877_),
    .A2(net57),
    .Z(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12962_ (.A1(_04875_),
    .A2(_04898_),
    .B(_04966_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12963_ (.A1(_04319_),
    .A2(_04789_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12964_ (.A1(_04894_),
    .A2(_04895_),
    .Z(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12965_ (.A1(_04894_),
    .A2(_04895_),
    .Z(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12966_ (.A1(_04890_),
    .A2(_04969_),
    .B(_04970_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12967_ (.I(_04889_),
    .Z(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12968_ (.I(_04972_),
    .Z(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12969_ (.A1(_04239_),
    .A2(_04973_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12970_ (.A1(_04968_),
    .A2(_04971_),
    .A3(_04974_),
    .Z(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12971_ (.A1(_04967_),
    .A2(_04975_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _12972_ (.A1(_04976_),
    .A2(_04965_),
    .ZN(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12973_ (.A1(_04962_),
    .A2(_04977_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _12974_ (.A1(_04808_),
    .A2(_04904_),
    .A3(_04978_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12975_ (.A1(_04500_),
    .A2(_04509_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12976_ (.I(_04519_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12977_ (.A1(_04500_),
    .A2(_04509_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12978_ (.A1(_04980_),
    .A2(_04981_),
    .B(_04982_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12979_ (.A1(_04484_),
    .A2(_04488_),
    .Z(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12980_ (.A1(_04730_),
    .A2(_04736_),
    .A3(_04745_),
    .Z(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12981_ (.A1(_04984_),
    .A2(_04985_),
    .Z(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12982_ (.A1(_04984_),
    .A2(_04985_),
    .Z(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _12983_ (.A1(_04983_),
    .A2(_04986_),
    .B(_04987_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12984_ (.A1(_04235_),
    .A2(_04799_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _12985_ (.A1(_04802_),
    .A2(_04989_),
    .A3(_04794_),
    .Z(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12986_ (.I(_04990_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12987_ (.A1(_04538_),
    .A2(_04447_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12988_ (.A1(_04512_),
    .A2(_04518_),
    .Z(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12989_ (.A1(_04512_),
    .A2(_04518_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12990_ (.A1(_04510_),
    .A2(_04993_),
    .B(_04994_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12991_ (.A1(_04648_),
    .A2(_04793_),
    .B(_04995_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12992_ (.A1(_04648_),
    .A2(_04793_),
    .A3(_04995_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12993_ (.A1(_04992_),
    .A2(_04996_),
    .B(_04997_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12994_ (.A1(_04991_),
    .A2(_04988_),
    .Z(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12995_ (.A1(_04998_),
    .A2(_04999_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _12996_ (.A1(_04988_),
    .A2(_04991_),
    .B(_05000_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12997_ (.A1(_04476_),
    .A2(_04489_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12998_ (.A1(_04839_),
    .A2(_04840_),
    .Z(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _12999_ (.A1(_05002_),
    .A2(_05003_),
    .Z(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13000_ (.A1(_04984_),
    .A2(_04983_),
    .A3(_04985_),
    .Z(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13001_ (.A1(_05002_),
    .A2(_05003_),
    .Z(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13002_ (.A1(_05004_),
    .A2(_05005_),
    .B(_05006_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13003_ (.A1(_04843_),
    .A2(_04842_),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13004_ (.A1(_05008_),
    .A2(_05007_),
    .Z(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13005_ (.A1(_04998_),
    .A2(_04999_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13006_ (.A1(_05004_),
    .A2(_05005_),
    .Z(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13007_ (.A1(_05006_),
    .A2(_05011_),
    .B(_05008_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13008_ (.A1(_05009_),
    .A2(_05010_),
    .B(_05012_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13009_ (.A1(_04845_),
    .A2(_04900_),
    .A3(_04902_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13010_ (.A1(_05013_),
    .A2(_05014_),
    .Z(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13011_ (.A1(_05013_),
    .A2(_05014_),
    .Z(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13012_ (.A1(_05001_),
    .A2(_05015_),
    .B(_05016_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13013_ (.A1(_04979_),
    .A2(_05017_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13014_ (.A1(_05001_),
    .A2(_05015_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13015_ (.A1(_04538_),
    .A2(_04672_),
    .A3(_04535_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13016_ (.A1(_04529_),
    .A2(_04540_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13017_ (.A1(_05020_),
    .A2(_05021_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13018_ (.A1(_04494_),
    .A2(_04520_),
    .Z(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13019_ (.A1(_04493_),
    .A2(_04521_),
    .B(_05023_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13020_ (.A1(_04795_),
    .A2(_04793_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13021_ (.A1(_04995_),
    .A2(_05025_),
    .A3(_04992_),
    .Z(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13022_ (.A1(_05024_),
    .A2(_05026_),
    .Z(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13023_ (.I(_05024_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13024_ (.A1(_05028_),
    .A2(_05026_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13025_ (.A1(_05022_),
    .A2(_05027_),
    .B(_05029_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13026_ (.I(_05030_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13027_ (.A1(_04493_),
    .A2(_04521_),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13028_ (.A1(_05005_),
    .A2(_05004_),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13029_ (.A1(_04490_),
    .A2(_05032_),
    .B(_05033_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13030_ (.A1(_05022_),
    .A2(_05027_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13031_ (.A1(_04490_),
    .A2(_05032_),
    .A3(_05033_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13032_ (.A1(_05034_),
    .A2(_05035_),
    .B(_05036_),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13033_ (.A1(_05010_),
    .A2(_05009_),
    .Z(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13034_ (.A1(_05037_),
    .A2(_05038_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13035_ (.A1(_05037_),
    .A2(_05038_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13036_ (.A1(_05031_),
    .A2(_05039_),
    .B(_05040_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13037_ (.A1(_05019_),
    .A2(_05041_),
    .Z(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13038_ (.A1(_05037_),
    .A2(_05038_),
    .A3(_05030_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13039_ (.I(_04523_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13040_ (.A1(_04523_),
    .A2(_04541_),
    .Z(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13041_ (.A1(_04528_),
    .A2(_05045_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13042_ (.A1(_05044_),
    .A2(_04541_),
    .B(_05046_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13043_ (.A1(_04410_),
    .A2(_04466_),
    .B(_04522_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _13044_ (.A1(_04410_),
    .A2(_04466_),
    .A3(_04522_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13045_ (.A1(_05048_),
    .A2(_04542_),
    .B(_05049_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13046_ (.A1(_04490_),
    .A2(_05032_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13047_ (.A1(_05022_),
    .A2(_05024_),
    .A3(_05026_),
    .Z(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13048_ (.A1(_05051_),
    .A2(_05033_),
    .A3(_05052_),
    .Z(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13049_ (.A1(_05050_),
    .A2(_05053_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13050_ (.A1(_05050_),
    .A2(_05053_),
    .Z(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13051_ (.A1(_05047_),
    .A2(_05054_),
    .B(_05055_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13052_ (.A1(_05056_),
    .A2(_05043_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13053_ (.A1(_05047_),
    .A2(_05054_),
    .Z(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13054_ (.A1(_04465_),
    .A2(_04543_),
    .Z(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13055_ (.A1(_04462_),
    .A2(_04544_),
    .B(_05059_),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13056_ (.A1(_05058_),
    .A2(_05060_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13057_ (.A1(_05061_),
    .A2(_05057_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _13058_ (.A1(_04723_),
    .A2(_05018_),
    .A3(_05042_),
    .A4(_05062_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13059_ (.A1(_05047_),
    .A2(_05054_),
    .Z(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13060_ (.A1(_05055_),
    .A2(_05064_),
    .B(_05043_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13061_ (.A1(_05058_),
    .A2(_05060_),
    .Z(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13062_ (.A1(_05043_),
    .A2(_05055_),
    .A3(_05064_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13063_ (.A1(_05065_),
    .A2(_05066_),
    .B(_05067_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _13064_ (.A1(_05018_),
    .A2(_05042_),
    .A3(_05068_),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13065_ (.A1(_04979_),
    .A2(_05017_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13066_ (.A1(_05037_),
    .A2(_05038_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13067_ (.A1(_05040_),
    .A2(_05030_),
    .A3(_05071_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13068_ (.A1(_04979_),
    .A2(_05017_),
    .B1(_05040_),
    .B2(_05072_),
    .C(_05019_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _13069_ (.A1(_05070_),
    .A2(_05073_),
    .Z(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13070_ (.I(_04892_),
    .Z(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13071_ (.I(_05075_),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13072_ (.I(_05076_),
    .Z(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13073_ (.A1(_04956_),
    .A2(_04957_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13074_ (.A1(_04956_),
    .A2(_04957_),
    .Z(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13075_ (.A1(_04953_),
    .A2(_05078_),
    .B(_05079_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13076_ (.A1(_04673_),
    .A2(_05077_),
    .A3(_05080_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13077_ (.I(_04973_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13078_ (.A1(_04671_),
    .A2(_05077_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13079_ (.A1(_05080_),
    .A2(_05083_),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13080_ (.A1(_04658_),
    .A2(_05082_),
    .A3(_05084_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13081_ (.A1(_05081_),
    .A2(_05085_),
    .Z(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13082_ (.A1(_04946_),
    .A2(_04950_),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13083_ (.A1(_04951_),
    .A2(_04958_),
    .B(_05087_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13084_ (.A1(_04929_),
    .A2(_04934_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13085_ (.A1(_04929_),
    .A2(_04934_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13086_ (.A1(_04924_),
    .A2(_05089_),
    .B(_05090_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13087_ (.A1(_04728_),
    .A2(_04305_),
    .B1(_04537_),
    .B2(_04266_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13088_ (.A1(_04728_),
    .A2(_04266_),
    .A3(_04305_),
    .A4(_04537_),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13089_ (.A1(_04947_),
    .A2(_05092_),
    .B(_05093_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13090_ (.A1(_04734_),
    .A2(_04781_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13091_ (.A1(_03400_),
    .A2(_04365_),
    .A3(_04431_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13092_ (.I(net48),
    .Z(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13093_ (.A1(_03384_),
    .A2(_05097_),
    .A3(_04371_),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13094_ (.A1(_05096_),
    .A2(_05098_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13095_ (.A1(_05095_),
    .A2(_05099_),
    .Z(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13096_ (.A1(_05094_),
    .A2(_05100_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13097_ (.I(_04954_),
    .Z(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13098_ (.I(_05102_),
    .Z(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13099_ (.A1(_04203_),
    .A2(_05103_),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13100_ (.I0(\filters.high[16] ),
    .I1(\filters.band[16] ),
    .S(_03189_),
    .Z(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13101_ (.I(_05105_),
    .Z(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _13102_ (.I(_05106_),
    .Z(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13103_ (.A1(_04513_),
    .A2(_05107_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13104_ (.A1(_04228_),
    .A2(_04788_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13105_ (.A1(_05104_),
    .A2(_05108_),
    .A3(_05109_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13106_ (.A1(_05101_),
    .A2(_05110_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13107_ (.A1(_05091_),
    .A2(_05111_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13108_ (.A1(_05091_),
    .A2(_05111_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13109_ (.A1(_05088_),
    .A2(_05112_),
    .B(_05113_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13110_ (.A1(_04320_),
    .A2(_05077_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13111_ (.A1(_05108_),
    .A2(_05109_),
    .Z(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13112_ (.A1(_05108_),
    .A2(_05109_),
    .Z(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13113_ (.A1(_05104_),
    .A2(_05116_),
    .B(_05117_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13114_ (.I(_05102_),
    .Z(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13115_ (.I(_05119_),
    .Z(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13116_ (.A1(_04796_),
    .A2(_05120_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13117_ (.A1(_05115_),
    .A2(_05118_),
    .A3(_05121_),
    .Z(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13118_ (.I(_05122_),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13119_ (.A1(_05114_),
    .A2(_05123_),
    .Z(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13120_ (.A1(_05114_),
    .A2(_05123_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13121_ (.A1(_05086_),
    .A2(_05124_),
    .B(_05125_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13122_ (.A1(_04908_),
    .A2(_04921_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13123_ (.A1(_04908_),
    .A2(_04921_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13124_ (.A1(_05127_),
    .A2(_04935_),
    .B(_05128_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13125_ (.A1(_04916_),
    .A2(_04920_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13126_ (.A1(_04913_),
    .A2(_04915_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13127_ (.A1(_03272_),
    .A2(_04273_),
    .A3(_04847_),
    .Z(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13128_ (.A1(_03254_),
    .A2(_04254_),
    .A3(_04910_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13129_ (.A1(\filters.cutoff_lut[16] ),
    .A2(_04468_),
    .Z(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13130_ (.I(_05134_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13131_ (.A1(_03201_),
    .A2(_04244_),
    .A3(_05135_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13132_ (.A1(_05132_),
    .A2(_05133_),
    .A3(_05136_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13133_ (.A1(_03317_),
    .A2(_04191_),
    .A3(_04470_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13134_ (.A1(net69),
    .A2(_04223_),
    .A3(_04812_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13135_ (.A1(_03303_),
    .A2(_04361_),
    .A3(_04816_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13136_ (.A1(_05138_),
    .A2(_05139_),
    .A3(_05140_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13137_ (.A1(_05131_),
    .A2(_05137_),
    .A3(_05141_),
    .Z(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13138_ (.A1(_05130_),
    .A2(_05142_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13139_ (.A1(_04931_),
    .A2(_04932_),
    .Z(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13140_ (.A1(_04930_),
    .A2(_04933_),
    .B(_05144_),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13141_ (.A1(_04362_),
    .A2(_04925_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13142_ (.A1(_04918_),
    .A2(_04919_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13143_ (.A1(_04918_),
    .A2(_04919_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13144_ (.A1(_05146_),
    .A2(_05147_),
    .B(_05148_),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13145_ (.I(_04397_),
    .Z(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13146_ (.A1(_05150_),
    .A2(_04304_),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13147_ (.A1(_03351_),
    .A2(_04751_),
    .A3(_04218_),
    .ZN(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13148_ (.A1(_03334_),
    .A2(net59),
    .A3(_04478_),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13149_ (.A1(_05152_),
    .A2(_05153_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13150_ (.A1(_05151_),
    .A2(_05154_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13151_ (.A1(_05145_),
    .A2(_05149_),
    .A3(_05155_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13152_ (.A1(_05143_),
    .A2(_05156_),
    .Z(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13153_ (.A1(_05129_),
    .A2(_05157_),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13154_ (.A1(_05088_),
    .A2(_05091_),
    .A3(_05111_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13155_ (.A1(_05129_),
    .A2(_05157_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13156_ (.A1(_05158_),
    .A2(_05159_),
    .B(_05160_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13157_ (.A1(_05130_),
    .A2(_05142_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13158_ (.A1(_05143_),
    .A2(_05156_),
    .B(_05162_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13159_ (.A1(_05131_),
    .A2(_05137_),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13160_ (.I(_05141_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13161_ (.A1(_05131_),
    .A2(_05137_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _13162_ (.A1(_05164_),
    .A2(_05165_),
    .B(_05166_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13163_ (.A1(_04400_),
    .A2(_04849_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13164_ (.A1(_05133_),
    .A2(_05136_),
    .Z(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13165_ (.A1(_05133_),
    .A2(_05136_),
    .Z(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _13166_ (.A1(_05168_),
    .A2(_05169_),
    .B(_05170_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13167_ (.A1(_04418_),
    .A2(_04848_),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13168_ (.A1(_04399_),
    .A2(_04911_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13169_ (.I(_05135_),
    .Z(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13170_ (.A1(_04349_),
    .A2(_05174_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _13171_ (.A1(_05172_),
    .A2(_05173_),
    .A3(_05175_),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13172_ (.A1(_04207_),
    .A2(_04471_),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13173_ (.A1(_04504_),
    .A2(_04813_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13174_ (.A1(_04415_),
    .A2(_04825_),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13175_ (.A1(_05177_),
    .A2(_05178_),
    .A3(_05179_),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13176_ (.A1(_05171_),
    .A2(_05176_),
    .A3(net41),
    .Z(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13177_ (.A1(_05152_),
    .A2(_05153_),
    .Z(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13178_ (.A1(_05151_),
    .A2(_05154_),
    .B(_05182_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13179_ (.A1(_05139_),
    .A2(_05140_),
    .Z(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13180_ (.A1(_05139_),
    .A2(_05140_),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _13181_ (.A1(_04193_),
    .A2(_04925_),
    .A3(_05184_),
    .B(_05185_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13182_ (.A1(_04353_),
    .A2(_04536_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13183_ (.A1(_03350_),
    .A2(_04218_),
    .A3(_04404_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13184_ (.A1(_03365_),
    .A2(_04751_),
    .A3(net53),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13185_ (.A1(_05188_),
    .A2(_05189_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13186_ (.A1(_05187_),
    .A2(_05190_),
    .Z(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13187_ (.A1(_05183_),
    .A2(_05186_),
    .A3(_05191_),
    .Z(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13188_ (.A1(_05167_),
    .A2(_05181_),
    .A3(_05192_),
    .Z(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13189_ (.A1(_05163_),
    .A2(_05193_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13190_ (.A1(_05094_),
    .A2(_05100_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13191_ (.A1(_05101_),
    .A2(_05110_),
    .B(_05195_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13192_ (.A1(_05149_),
    .A2(_05155_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13193_ (.A1(_05149_),
    .A2(_05155_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13194_ (.A1(_05145_),
    .A2(_05197_),
    .B(_05198_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13195_ (.A1(_05096_),
    .A2(_05098_),
    .Z(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13196_ (.A1(_05095_),
    .A2(_05099_),
    .B(_05200_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13197_ (.A1(_04258_),
    .A2(_04768_),
    .ZN(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13198_ (.A1(_05097_),
    .A2(_04432_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13199_ (.A1(_04732_),
    .A2(_04516_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13200_ (.A1(_05202_),
    .A2(_05203_),
    .A3(_05204_),
    .Z(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13201_ (.A1(_05201_),
    .A2(_05205_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13202_ (.I(_03189_),
    .Z(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13203_ (.A1(\filters.band[16] ),
    .A2(_05207_),
    .Z(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13204_ (.A1(\filters.high[16] ),
    .A2(_03472_),
    .B(_05208_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13205_ (.A1(_04562_),
    .A2(_05209_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13206_ (.I(_04225_),
    .Z(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13207_ (.I(_04771_),
    .Z(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13208_ (.A1(_05211_),
    .A2(_05212_),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13209_ (.I0(\filters.high[17] ),
    .I1(\filters.band[17] ),
    .S(_03188_),
    .Z(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13210_ (.I(_05214_),
    .Z(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13211_ (.I(_05215_),
    .Z(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13212_ (.A1(_04307_),
    .A2(_05216_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13213_ (.A1(_05210_),
    .A2(_05213_),
    .A3(_05217_),
    .Z(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13214_ (.A1(_05206_),
    .A2(_05218_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13215_ (.A1(_05196_),
    .A2(_05199_),
    .A3(_05219_),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13216_ (.A1(_05194_),
    .A2(_05220_),
    .Z(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13217_ (.A1(_05161_),
    .A2(net52),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13218_ (.A1(_05086_),
    .A2(_05114_),
    .A3(_05123_),
    .Z(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13219_ (.A1(_05161_),
    .A2(net52),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13220_ (.A1(_05222_),
    .A2(_05223_),
    .B(_05224_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13221_ (.A1(_05163_),
    .A2(_05193_),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13222_ (.A1(_05194_),
    .A2(_05220_),
    .B(_05226_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13223_ (.A1(_05167_),
    .A2(_05181_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13224_ (.I(_05183_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13225_ (.A1(_05229_),
    .A2(_05186_),
    .A3(_05191_),
    .Z(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13226_ (.A1(_05167_),
    .A2(_05181_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13227_ (.A1(_05228_),
    .A2(_05230_),
    .B(_05231_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13228_ (.A1(_05171_),
    .A2(_05176_),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13229_ (.I(_05180_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13230_ (.A1(_05171_),
    .A2(_05176_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13231_ (.A1(_05233_),
    .A2(_05234_),
    .B(_05235_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13232_ (.A1(_04400_),
    .A2(_04912_),
    .B1(_05174_),
    .B2(_04349_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13233_ (.A1(_04349_),
    .A2(_04399_),
    .A3(_04912_),
    .A4(_05174_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13234_ (.A1(_05172_),
    .A2(_05237_),
    .B(_05238_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13235_ (.A1(_04310_),
    .A2(_04848_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13236_ (.A1(_03287_),
    .A2(_04222_),
    .A3(_04910_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13237_ (.A1(_03272_),
    .A2(_04273_),
    .A3(_05134_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13238_ (.A1(_05241_),
    .A2(_05242_),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13239_ (.A1(_05240_),
    .A2(_05243_),
    .Z(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13240_ (.A1(_05239_),
    .A2(_05244_),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13241_ (.A1(_04511_),
    .A2(_04824_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _13242_ (.A1(net43),
    .A2(_04208_),
    .A3(_04855_),
    .A4(_04825_),
    .Z(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _13243_ (.A1(net44),
    .A2(_04855_),
    .B1(_04825_),
    .B2(_04208_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _13244_ (.A1(_05246_),
    .A2(_05247_),
    .A3(_05248_),
    .Z(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13245_ (.A1(_05247_),
    .A2(_05248_),
    .B(_05246_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13246_ (.A1(_05249_),
    .A2(_05250_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13247_ (.A1(_05245_),
    .A2(_05251_),
    .Z(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13248_ (.A1(_05188_),
    .A2(_05189_),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13249_ (.A1(_05187_),
    .A2(_05190_),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13250_ (.A1(_05254_),
    .A2(_05253_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13251_ (.I(_04817_),
    .Z(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13252_ (.I(_04414_),
    .Z(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13253_ (.A1(_04422_),
    .A2(_04856_),
    .B1(_05256_),
    .B2(_05257_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13254_ (.A1(_04311_),
    .A2(_05257_),
    .A3(_04856_),
    .A4(_05256_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13255_ (.A1(_05177_),
    .A2(_05258_),
    .B(_05259_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13256_ (.I(_04432_),
    .Z(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13257_ (.A1(_04353_),
    .A2(_05261_),
    .Z(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13258_ (.A1(_03365_),
    .A2(net53),
    .A3(_04478_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13259_ (.A1(_03384_),
    .A2(_04344_),
    .A3(_04372_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13260_ (.A1(_05263_),
    .A2(_05264_),
    .Z(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13261_ (.A1(_05262_),
    .A2(_05265_),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13262_ (.A1(_05255_),
    .A2(_05260_),
    .A3(_05266_),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13263_ (.A1(_05236_),
    .A2(_05252_),
    .A3(_05267_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13264_ (.A1(_05095_),
    .A2(_05099_),
    .Z(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13265_ (.A1(_05200_),
    .A2(_05269_),
    .B(_05205_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13266_ (.A1(_05206_),
    .A2(_05218_),
    .B(_05270_),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13267_ (.A1(_05186_),
    .A2(_05191_),
    .ZN(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13268_ (.A1(_05186_),
    .A2(_05191_),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13269_ (.A1(_05229_),
    .A2(_05272_),
    .B(_05273_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13270_ (.A1(_04288_),
    .A2(_05261_),
    .B1(_04517_),
    .B2(_04421_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13271_ (.A1(_04288_),
    .A2(_04421_),
    .A3(_05261_),
    .A4(_04781_),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13272_ (.A1(_05202_),
    .A2(_05275_),
    .B(_05276_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13273_ (.A1(_04258_),
    .A2(_04771_),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13274_ (.A1(_05097_),
    .A2(_04780_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13275_ (.A1(_04249_),
    .A2(_04741_),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13276_ (.A1(_05278_),
    .A2(_05279_),
    .A3(_05280_),
    .Z(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13277_ (.A1(_05277_),
    .A2(_05281_),
    .ZN(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13278_ (.A1(_04296_),
    .A2(_05216_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13279_ (.A1(_04226_),
    .A2(_04893_),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13280_ (.I0(\filters.high[18] ),
    .I1(\filters.band[18] ),
    .S(_03188_),
    .Z(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13281_ (.I(_05285_),
    .Z(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13282_ (.A1(_04373_),
    .A2(_05286_),
    .ZN(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13283_ (.A1(_05284_),
    .A2(_05287_),
    .Z(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13284_ (.A1(_05283_),
    .A2(_05288_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13285_ (.A1(_05282_),
    .A2(_05289_),
    .Z(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13286_ (.A1(_05271_),
    .A2(_05274_),
    .A3(_05290_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13287_ (.A1(_05232_),
    .A2(_05268_),
    .A3(_05291_),
    .Z(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13288_ (.A1(_05292_),
    .A2(_05227_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13289_ (.I(_05120_),
    .Z(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13290_ (.A1(_04797_),
    .A2(_05294_),
    .B(_05118_),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13291_ (.A1(_04797_),
    .A2(_05294_),
    .A3(_05118_),
    .ZN(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13292_ (.A1(_05115_),
    .A2(_05295_),
    .B(_05296_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13293_ (.A1(_05199_),
    .A2(_05219_),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13294_ (.A1(_05199_),
    .A2(_05219_),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13295_ (.A1(net46),
    .A2(_05298_),
    .B(_05299_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13296_ (.A1(_04586_),
    .A2(_05294_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13297_ (.A1(_05213_),
    .A2(_05217_),
    .ZN(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13298_ (.A1(_05213_),
    .A2(_05217_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13299_ (.A1(_05210_),
    .A2(_05302_),
    .B(_05303_),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13300_ (.I(_05106_),
    .Z(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13301_ (.I(_05305_),
    .Z(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13302_ (.I(_05306_),
    .Z(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13303_ (.A1(_04238_),
    .A2(_05307_),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13304_ (.A1(_05304_),
    .A2(_05308_),
    .Z(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13305_ (.A1(_05301_),
    .A2(_05309_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13306_ (.A1(_05297_),
    .A2(_05300_),
    .A3(_05310_),
    .Z(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13307_ (.A1(_05311_),
    .A2(_05293_),
    .Z(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13308_ (.A1(_05312_),
    .A2(_05225_),
    .Z(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13309_ (.A1(_05225_),
    .A2(_05312_),
    .Z(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13310_ (.A1(_05126_),
    .A2(net40),
    .B(_05314_),
    .ZN(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13311_ (.I(_05310_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13312_ (.A1(_05300_),
    .A2(_05316_),
    .Z(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13313_ (.A1(_05297_),
    .A2(_05317_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13314_ (.A1(_05300_),
    .A2(_05316_),
    .B(_05318_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13315_ (.A1(_05227_),
    .A2(_05292_),
    .ZN(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13316_ (.A1(_05293_),
    .A2(_05311_),
    .B(_05320_),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13317_ (.A1(_05232_),
    .A2(_05268_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13318_ (.I(_05291_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13319_ (.A1(_05232_),
    .A2(_05268_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13320_ (.A1(_05322_),
    .A2(_05323_),
    .B(_05324_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13321_ (.A1(_05236_),
    .A2(_05252_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13322_ (.I(_05267_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13323_ (.A1(_05236_),
    .A2(_05252_),
    .ZN(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13324_ (.A1(_05326_),
    .A2(_05327_),
    .B(_05328_),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13325_ (.A1(_05239_),
    .A2(_05244_),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13326_ (.A1(_05245_),
    .A2(_05251_),
    .B(_05330_),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13327_ (.A1(_05241_),
    .A2(_05242_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13328_ (.A1(_05240_),
    .A2(_05243_),
    .B(_05332_),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13329_ (.A1(_04413_),
    .A2(_04847_),
    .ZN(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13330_ (.A1(_03302_),
    .A2(_04309_),
    .A3(_04909_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13331_ (.A1(_03287_),
    .A2(_04221_),
    .A3(_05134_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13332_ (.A1(_05335_),
    .A2(_05336_),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13333_ (.A1(_05334_),
    .A2(_05337_),
    .Z(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13334_ (.A1(_05333_),
    .A2(_05338_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13335_ (.A1(_04302_),
    .A2(_04471_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _13336_ (.A1(_04297_),
    .A2(_04207_),
    .A3(_04814_),
    .A4(_04834_),
    .Z(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _13337_ (.A1(_04502_),
    .A2(_04814_),
    .B1(_04817_),
    .B2(_04297_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _13338_ (.A1(_05340_),
    .A2(_05341_),
    .A3(_05342_),
    .Z(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13339_ (.A1(_05341_),
    .A2(_05342_),
    .B(_05340_),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13340_ (.A1(_05343_),
    .A2(_05344_),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13341_ (.A1(_05345_),
    .A2(_05339_),
    .Z(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13342_ (.A1(_05346_),
    .A2(_05331_),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13343_ (.A1(_05262_),
    .A2(_05265_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13344_ (.A1(_05263_),
    .A2(_05264_),
    .B(_05348_),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13345_ (.I(_04813_),
    .Z(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _13346_ (.A1(_04725_),
    .A2(_04760_),
    .A3(_05350_),
    .A4(_04835_),
    .ZN(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13347_ (.A1(_05246_),
    .A2(_05248_),
    .B(_05351_),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13348_ (.A1(_04352_),
    .A2(_04515_),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13349_ (.A1(_04425_),
    .A2(_04404_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13350_ (.A1(_04751_),
    .A2(_04432_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13351_ (.A1(_05353_),
    .A2(_05354_),
    .A3(_05355_),
    .Z(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13352_ (.A1(_05356_),
    .A2(_05352_),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13353_ (.A1(_05349_),
    .A2(_05357_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13354_ (.A1(_05358_),
    .A2(_05347_),
    .Z(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13355_ (.I(_05277_),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13356_ (.A1(_05282_),
    .A2(_05289_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13357_ (.A1(_05360_),
    .A2(_05281_),
    .B(_05361_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13358_ (.A1(_05260_),
    .A2(_05266_),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13359_ (.A1(_05260_),
    .A2(_05266_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13360_ (.A1(net64),
    .A2(_05363_),
    .B(_05364_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13361_ (.A1(_04417_),
    .A2(_04516_),
    .B1(_04741_),
    .B2(_04732_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13362_ (.A1(_04287_),
    .A2(_04249_),
    .A3(_04516_),
    .A4(_04741_),
    .ZN(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13363_ (.A1(_05278_),
    .A2(_05366_),
    .B(_05367_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13364_ (.A1(net63),
    .A2(_04891_),
    .ZN(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13365_ (.A1(net49),
    .A2(_04740_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13366_ (.A1(_04248_),
    .A2(_04770_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13367_ (.A1(_05369_),
    .A2(_05370_),
    .A3(_05371_),
    .Z(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13368_ (.A1(_05372_),
    .A2(_05368_),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13369_ (.I(_05285_),
    .Z(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13370_ (.A1(_04295_),
    .A2(_05374_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13371_ (.A1(_04225_),
    .A2(_04954_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13372_ (.I0(\filters.high[19] ),
    .I1(\filters.band[19] ),
    .S(_04739_),
    .Z(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13373_ (.I(_05377_),
    .Z(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13374_ (.A1(_04213_),
    .A2(_05378_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13375_ (.A1(_05376_),
    .A2(_05379_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13376_ (.A1(_05375_),
    .A2(_05380_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13377_ (.A1(_05381_),
    .A2(_05373_),
    .Z(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13378_ (.A1(_05382_),
    .A2(_05365_),
    .Z(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13379_ (.A1(_05383_),
    .A2(_05362_),
    .Z(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13380_ (.A1(_05329_),
    .A2(_05359_),
    .A3(_05384_),
    .Z(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13381_ (.A1(_04526_),
    .A2(_05120_),
    .A3(_05309_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13382_ (.A1(_05304_),
    .A2(_05308_),
    .B(_05386_),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13383_ (.I(_05271_),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13384_ (.A1(_05274_),
    .A2(_05290_),
    .Z(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13385_ (.A1(_05274_),
    .A2(_05290_),
    .Z(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13386_ (.A1(_05388_),
    .A2(_05389_),
    .B(_05390_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13387_ (.A1(_04526_),
    .A2(_05307_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13388_ (.A1(_05284_),
    .A2(_05287_),
    .Z(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13389_ (.I(_05214_),
    .Z(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13390_ (.I(_05394_),
    .Z(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13391_ (.I(_05395_),
    .Z(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13392_ (.A1(_04624_),
    .A2(_05396_),
    .A3(_05288_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13393_ (.A1(_05393_),
    .A2(_05397_),
    .Z(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13394_ (.I(_05396_),
    .Z(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13395_ (.A1(_04671_),
    .A2(_05399_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13396_ (.A1(_05398_),
    .A2(_05400_),
    .Z(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13397_ (.A1(_05392_),
    .A2(_05401_),
    .Z(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13398_ (.A1(_05387_),
    .A2(_05391_),
    .A3(_05402_),
    .Z(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13399_ (.A1(_05325_),
    .A2(_05385_),
    .A3(_05403_),
    .ZN(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13400_ (.A1(_05404_),
    .A2(_05321_),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13401_ (.A1(_05405_),
    .A2(_05319_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13402_ (.A1(_05406_),
    .A2(_05315_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13403_ (.A1(_05313_),
    .A2(_05126_),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13404_ (.A1(_04943_),
    .A2(_04959_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13405_ (.A1(_04943_),
    .A2(_04959_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13406_ (.A1(_04940_),
    .A2(_05409_),
    .B(_05410_),
    .ZN(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13407_ (.A1(_04658_),
    .A2(_05082_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13408_ (.A1(_05412_),
    .A2(_05084_),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13409_ (.I(_05413_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13410_ (.A1(_04673_),
    .A2(_05082_),
    .B(_04971_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13411_ (.A1(_04673_),
    .A2(_05082_),
    .A3(_04971_),
    .ZN(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13412_ (.A1(_04968_),
    .A2(_05415_),
    .B(_05416_),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13413_ (.A1(_05411_),
    .A2(_05414_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13414_ (.A1(_05417_),
    .A2(_05418_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13415_ (.A1(_05411_),
    .A2(_05414_),
    .B(_05419_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13416_ (.A1(_04907_),
    .A2(_04936_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13417_ (.A1(_04907_),
    .A2(_04936_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13418_ (.A1(_05421_),
    .A2(_04960_),
    .B(_05422_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13419_ (.A1(_05158_),
    .A2(_05159_),
    .Z(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13420_ (.A1(_05423_),
    .A2(_05424_),
    .ZN(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13421_ (.A1(_05417_),
    .A2(_05411_),
    .A3(_05413_),
    .Z(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13422_ (.A1(_05423_),
    .A2(_05424_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13423_ (.A1(_05425_),
    .A2(_05426_),
    .B(_05427_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13424_ (.A1(_05161_),
    .A2(_05221_),
    .A3(_05223_),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13425_ (.A1(_05428_),
    .A2(_05429_),
    .Z(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13426_ (.A1(_05428_),
    .A2(net62),
    .Z(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13427_ (.A1(_05420_),
    .A2(_05430_),
    .B(_05431_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13428_ (.A1(_05432_),
    .A2(_05408_),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13429_ (.A1(_05420_),
    .A2(_05430_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13430_ (.I(_04967_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13431_ (.A1(_05435_),
    .A2(_04975_),
    .ZN(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13432_ (.A1(_04965_),
    .A2(_04976_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13433_ (.A1(_05436_),
    .A2(_05437_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13434_ (.A1(_04906_),
    .A2(_04961_),
    .Z(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13435_ (.A1(_04962_),
    .A2(_04977_),
    .B(_05439_),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13436_ (.A1(_05423_),
    .A2(_05424_),
    .A3(_05426_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13437_ (.A1(_05440_),
    .A2(_05441_),
    .Z(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13438_ (.A1(_05440_),
    .A2(_05441_),
    .Z(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13439_ (.A1(_05438_),
    .A2(_05442_),
    .B(_05443_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13440_ (.A1(_05434_),
    .A2(_05444_),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13441_ (.A1(_05442_),
    .A2(_05438_),
    .ZN(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13442_ (.A1(_04904_),
    .A2(_04978_),
    .Z(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13443_ (.A1(_04904_),
    .A2(_04978_),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13444_ (.A1(_04808_),
    .A2(_05447_),
    .B(_05448_),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13445_ (.A1(_05446_),
    .A2(_05449_),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _13446_ (.A1(_05407_),
    .A2(_05433_),
    .A3(_05445_),
    .A4(_05450_),
    .ZN(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _13447_ (.A1(_05063_),
    .A2(_05069_),
    .A3(_05074_),
    .B(_05451_),
    .ZN(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13448_ (.A1(_05315_),
    .A2(_05406_),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13449_ (.A1(_05408_),
    .A2(_05432_),
    .ZN(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13450_ (.A1(_05407_),
    .A2(_05433_),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13451_ (.A1(_05434_),
    .A2(_05444_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13452_ (.A1(_05434_),
    .A2(_05444_),
    .B1(_05446_),
    .B2(_05449_),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13453_ (.A1(_05456_),
    .A2(_05457_),
    .Z(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13454_ (.A1(_05315_),
    .A2(_05406_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _13455_ (.A1(_05453_),
    .A2(_05454_),
    .B1(_05455_),
    .B2(_05458_),
    .C(_05459_),
    .ZN(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _13456_ (.A1(_05452_),
    .A2(_05460_),
    .Z(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13457_ (.A1(_05391_),
    .A2(_05402_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13458_ (.A1(_05391_),
    .A2(_05402_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13459_ (.A1(_05387_),
    .A2(_05462_),
    .B(_05463_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13460_ (.A1(_05325_),
    .A2(_05385_),
    .ZN(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13461_ (.I(_05403_),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13462_ (.A1(_05325_),
    .A2(_05385_),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13463_ (.A1(_05465_),
    .A2(_05466_),
    .B(_05467_),
    .ZN(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13464_ (.A1(_04669_),
    .A2(_05307_),
    .A3(_05401_),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13465_ (.A1(_05398_),
    .A2(_05400_),
    .B(_05469_),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13466_ (.A1(_05365_),
    .A2(_05382_),
    .Z(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13467_ (.A1(_05362_),
    .A2(_05383_),
    .B(_05471_),
    .ZN(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13468_ (.A1(_04586_),
    .A2(_05399_),
    .ZN(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13469_ (.I(_05374_),
    .Z(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13470_ (.I(_05474_),
    .Z(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13471_ (.A1(_04625_),
    .A2(_05475_),
    .A3(_05380_),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13472_ (.A1(_05376_),
    .A2(_05379_),
    .B(_05476_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13473_ (.A1(_04672_),
    .A2(_05475_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13474_ (.A1(_05477_),
    .A2(_05478_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13475_ (.A1(_05473_),
    .A2(_05479_),
    .Z(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13476_ (.A1(_05472_),
    .A2(_05480_),
    .Z(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13477_ (.A1(_05470_),
    .A2(_05481_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13478_ (.A1(_05329_),
    .A2(_05359_),
    .Z(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13479_ (.A1(_05329_),
    .A2(_05359_),
    .Z(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13480_ (.A1(_05483_),
    .A2(_05384_),
    .B(_05484_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13481_ (.A1(_05331_),
    .A2(_05346_),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13482_ (.A1(_05347_),
    .A2(_05358_),
    .B(_05486_),
    .ZN(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13483_ (.A1(_05354_),
    .A2(_05355_),
    .Z(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13484_ (.A1(_05354_),
    .A2(_05355_),
    .Z(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13485_ (.A1(_05353_),
    .A2(_05488_),
    .B(_05489_),
    .ZN(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13486_ (.I(_05350_),
    .Z(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13487_ (.I(_05491_),
    .Z(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13488_ (.I(_05256_),
    .Z(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _13489_ (.A1(_04299_),
    .A2(_04210_),
    .A3(_05492_),
    .A4(_05493_),
    .ZN(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13490_ (.A1(_05340_),
    .A2(_05342_),
    .B(_05494_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13491_ (.I(_04768_),
    .Z(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13492_ (.A1(_05150_),
    .A2(_05496_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13493_ (.A1(_04479_),
    .A2(_05261_),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13494_ (.I(_04752_),
    .Z(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13495_ (.A1(_05499_),
    .A2(_04782_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13496_ (.A1(_05497_),
    .A2(_05498_),
    .A3(_05500_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13497_ (.A1(_05495_),
    .A2(_05501_),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13498_ (.A1(_05502_),
    .A2(_05490_),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13499_ (.A1(_05333_),
    .A2(_05338_),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13500_ (.A1(_05339_),
    .A2(_05345_),
    .B(_05504_),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13501_ (.A1(_04537_),
    .A2(_04472_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13502_ (.A1(_03352_),
    .A2(_04219_),
    .A3(_05350_),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13503_ (.A1(_03366_),
    .A2(_04885_),
    .A3(_04835_),
    .ZN(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13504_ (.A1(_05507_),
    .A2(_05508_),
    .Z(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13505_ (.A1(_05506_),
    .A2(_05509_),
    .Z(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13506_ (.A1(_05335_),
    .A2(_05336_),
    .Z(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13507_ (.A1(_05334_),
    .A2(_05337_),
    .B(_05511_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13508_ (.A1(_04502_),
    .A2(_04914_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13509_ (.I(_05135_),
    .Z(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13510_ (.A1(_04504_),
    .A2(_05514_),
    .ZN(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13511_ (.I(_04912_),
    .Z(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13512_ (.A1(_04507_),
    .A2(_05516_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13513_ (.A1(_05513_),
    .A2(_05515_),
    .A3(_05517_),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13514_ (.A1(_05512_),
    .A2(_05518_),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13515_ (.A1(_05510_),
    .A2(_05519_),
    .Z(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13516_ (.A1(_05505_),
    .A2(_05520_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13517_ (.A1(_05503_),
    .A2(_05521_),
    .Z(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13518_ (.A1(_05487_),
    .A2(_05522_),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13519_ (.I(_05368_),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13520_ (.A1(_05524_),
    .A2(_05372_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13521_ (.A1(net45),
    .A2(_05381_),
    .B(_05525_),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13522_ (.A1(_05351_),
    .A2(_05249_),
    .B(_05356_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13523_ (.A1(_05349_),
    .A2(net61),
    .B(_05527_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13524_ (.I(_05378_),
    .Z(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13525_ (.I(_05529_),
    .Z(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13526_ (.A1(_04551_),
    .A2(_05530_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13527_ (.A1(_04326_),
    .A2(_05107_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13528_ (.I0(\filters.high[20] ),
    .I1(\filters.band[20] ),
    .S(_03189_),
    .Z(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13529_ (.I(_05533_),
    .Z(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13530_ (.A1(_04307_),
    .A2(_05534_),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13531_ (.A1(_05532_),
    .A2(_05535_),
    .Z(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13532_ (.A1(_05531_),
    .A2(_05536_),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13533_ (.I(_04495_),
    .Z(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13534_ (.I(_04742_),
    .Z(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13535_ (.I(_04881_),
    .Z(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13536_ (.A1(_05538_),
    .A2(_05539_),
    .B1(_04973_),
    .B2(_05540_),
    .ZN(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13537_ (.A1(_05538_),
    .A2(_05540_),
    .A3(_05539_),
    .A4(_04973_),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13538_ (.A1(_05369_),
    .A2(_05541_),
    .B(_05542_),
    .ZN(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13539_ (.A1(_04734_),
    .A2(_05102_),
    .ZN(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13540_ (.A1(_04270_),
    .A2(_05212_),
    .ZN(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13541_ (.A1(_04881_),
    .A2(_04952_),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13542_ (.A1(_05544_),
    .A2(_05545_),
    .A3(_05546_),
    .Z(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13543_ (.A1(_05543_),
    .A2(_05547_),
    .ZN(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13544_ (.A1(_05537_),
    .A2(_05548_),
    .ZN(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13545_ (.A1(_05528_),
    .A2(_05549_),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13546_ (.A1(_05526_),
    .A2(_05550_),
    .Z(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13547_ (.A1(_05523_),
    .A2(_05551_),
    .Z(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _13548_ (.A1(_05482_),
    .A2(_05485_),
    .A3(_05552_),
    .Z(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _13549_ (.A1(_05464_),
    .A2(_05468_),
    .A3(_05553_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13550_ (.I(_05321_),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13551_ (.A1(_05319_),
    .A2(_05405_),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _13552_ (.A1(_05555_),
    .A2(net39),
    .B(_05556_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13553_ (.A1(_05554_),
    .A2(_05557_),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13554_ (.A1(_05461_),
    .A2(_05558_),
    .Z(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13555_ (.I(_05559_),
    .Z(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13556_ (.I(\filters.low[0] ),
    .Z(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13557_ (.A1(_05561_),
    .A2(_03348_),
    .ZN(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13558_ (.A1(\filters.band[0] ),
    .A2(_03473_),
    .ZN(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _13559_ (.A1(_05560_),
    .A2(_05562_),
    .A3(_05563_),
    .Z(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13560_ (.A1(_05562_),
    .A2(_05563_),
    .B(_05560_),
    .ZN(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13561_ (.A1(_05564_),
    .A2(_05565_),
    .ZN(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13562_ (.I(_04187_),
    .Z(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13563_ (.A1(\filters.band[0] ),
    .A2(_05567_),
    .B(_03753_),
    .ZN(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13564_ (.A1(_04189_),
    .A2(_05566_),
    .B(_05568_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13565_ (.A1(_03758_),
    .A2(_03479_),
    .ZN(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13566_ (.I(_05569_),
    .Z(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13567_ (.I(_05570_),
    .Z(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13568_ (.I(_05569_),
    .Z(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13569_ (.I(_05572_),
    .Z(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13570_ (.A1(_05560_),
    .A2(_05562_),
    .A3(_05563_),
    .ZN(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13571_ (.A1(_05554_),
    .A2(_05557_),
    .Z(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13572_ (.A1(net35),
    .A2(net36),
    .B(_05558_),
    .ZN(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13573_ (.A1(_05468_),
    .A2(_05553_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13574_ (.A1(_05468_),
    .A2(_05553_),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13575_ (.A1(_05464_),
    .A2(_05577_),
    .B(_05578_),
    .ZN(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13576_ (.A1(_05472_),
    .A2(_05480_),
    .ZN(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13577_ (.A1(_05470_),
    .A2(_05481_),
    .B(_05580_),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13578_ (.A1(_05523_),
    .A2(_05551_),
    .Z(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13579_ (.A1(_05523_),
    .A2(_05551_),
    .ZN(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13580_ (.A1(_05485_),
    .A2(_05552_),
    .Z(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _13581_ (.A1(_05485_),
    .A2(_05582_),
    .A3(_05583_),
    .B1(_05584_),
    .B2(_05482_),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13582_ (.I(_04675_),
    .Z(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13583_ (.I(_05475_),
    .Z(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13584_ (.A1(_05586_),
    .A2(_05587_),
    .A3(_05477_),
    .ZN(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13585_ (.I(_04587_),
    .Z(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13586_ (.A1(_05589_),
    .A2(_05399_),
    .A3(_05479_),
    .ZN(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13587_ (.A1(_05588_),
    .A2(_05590_),
    .Z(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13588_ (.A1(_05528_),
    .A2(_05549_),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13589_ (.A1(_05526_),
    .A2(_05550_),
    .ZN(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13590_ (.A1(_05592_),
    .A2(_05593_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13591_ (.A1(_04659_),
    .A2(_05587_),
    .ZN(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13592_ (.I(_05530_),
    .Z(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13593_ (.A1(_04644_),
    .A2(_05596_),
    .A3(_05536_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13594_ (.A1(_05532_),
    .A2(_05535_),
    .B(_05597_),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13595_ (.A1(_04796_),
    .A2(_05596_),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13596_ (.A1(_05598_),
    .A2(_05599_),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13597_ (.A1(_05595_),
    .A2(_05600_),
    .Z(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13598_ (.A1(_05594_),
    .A2(_05601_),
    .ZN(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13599_ (.A1(_05591_),
    .A2(_05602_),
    .Z(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13600_ (.A1(_05487_),
    .A2(_05522_),
    .Z(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13601_ (.A1(_05523_),
    .A2(_05551_),
    .B(_05604_),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13602_ (.I(_05543_),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13603_ (.A1(_05606_),
    .A2(_05547_),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13604_ (.A1(_05537_),
    .A2(_05548_),
    .B(_05607_),
    .ZN(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13605_ (.A1(_05494_),
    .A2(_05343_),
    .B(_05501_),
    .ZN(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13606_ (.A1(_05490_),
    .A2(_05502_),
    .B(_05609_),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13607_ (.A1(_04204_),
    .A2(_05534_),
    .ZN(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13608_ (.A1(_04325_),
    .A2(_05215_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13609_ (.I0(\filters.high[21] ),
    .I1(\filters.band[21] ),
    .S(_05207_),
    .Z(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13610_ (.A1(_04306_),
    .A2(_05613_),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13611_ (.A1(_05612_),
    .A2(_05614_),
    .Z(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13612_ (.A1(_05611_),
    .A2(_05615_),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13613_ (.I(_04889_),
    .Z(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13614_ (.A1(_04879_),
    .A2(_05617_),
    .B1(_04952_),
    .B2(_04878_),
    .ZN(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13615_ (.A1(_04879_),
    .A2(_04881_),
    .A3(_04972_),
    .A4(_05075_),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13616_ (.A1(_05544_),
    .A2(_05618_),
    .B(_05619_),
    .ZN(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13617_ (.A1(_04501_),
    .A2(_05105_),
    .Z(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13618_ (.A1(_04269_),
    .A2(_04892_),
    .Z(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13619_ (.A1(_04506_),
    .A2(_04954_),
    .Z(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13620_ (.A1(_05621_),
    .A2(_05622_),
    .A3(_05623_),
    .Z(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13621_ (.A1(_05620_),
    .A2(_05624_),
    .Z(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13622_ (.A1(_05616_),
    .A2(_05625_),
    .ZN(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13623_ (.A1(_05610_),
    .A2(_05626_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13624_ (.A1(_05608_),
    .A2(_05627_),
    .Z(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13625_ (.A1(_05505_),
    .A2(_05520_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13626_ (.A1(_05503_),
    .A2(_05521_),
    .B(_05629_),
    .ZN(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13627_ (.A1(_05498_),
    .A2(_05500_),
    .Z(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13628_ (.A1(_05498_),
    .A2(_05500_),
    .Z(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13629_ (.A1(_05497_),
    .A2(_05631_),
    .B(_05632_),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13630_ (.A1(_05507_),
    .A2(_05508_),
    .Z(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13631_ (.A1(_05507_),
    .A2(_05508_),
    .Z(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13632_ (.A1(_05506_),
    .A2(_05634_),
    .B(_05635_),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13633_ (.A1(_05150_),
    .A2(_05212_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13634_ (.A1(_04479_),
    .A2(_04781_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13635_ (.A1(_05499_),
    .A2(_04742_),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13636_ (.A1(_05637_),
    .A2(_05638_),
    .A3(_05639_),
    .Z(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13637_ (.A1(_05636_),
    .A2(_05640_),
    .ZN(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13638_ (.A1(_05633_),
    .A2(_05641_),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13639_ (.A1(_05512_),
    .A2(_05518_),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13640_ (.A1(_05510_),
    .A2(_05519_),
    .B(_05643_),
    .ZN(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13641_ (.A1(_04434_),
    .A2(_04473_),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13642_ (.A1(_03366_),
    .A2(_04885_),
    .A3(_05350_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13643_ (.A1(_03385_),
    .A2(_04372_),
    .A3(_04835_),
    .ZN(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13644_ (.A1(_05646_),
    .A2(_05647_),
    .Z(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13645_ (.A1(_05645_),
    .A2(_05648_),
    .Z(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13646_ (.I(_05516_),
    .Z(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13647_ (.I(_05174_),
    .Z(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13648_ (.I(_05651_),
    .Z(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13649_ (.A1(_05257_),
    .A2(_05650_),
    .B1(_05652_),
    .B2(_04422_),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13650_ (.I(_04911_),
    .Z(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13651_ (.I(_05654_),
    .Z(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13652_ (.I(_05514_),
    .Z(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13653_ (.A1(_04497_),
    .A2(_05257_),
    .A3(_05655_),
    .A4(_05656_),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13654_ (.A1(_05513_),
    .A2(_05653_),
    .B(_05657_),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13655_ (.A1(_04511_),
    .A2(_04914_),
    .ZN(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13656_ (.A1(_03318_),
    .A2(_04191_),
    .A3(_05514_),
    .ZN(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13657_ (.A1(_03334_),
    .A2(_04548_),
    .A3(_05516_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13658_ (.A1(_05659_),
    .A2(_05660_),
    .A3(_05661_),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13659_ (.A1(_05658_),
    .A2(_05662_),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13660_ (.A1(_05649_),
    .A2(_05663_),
    .Z(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13661_ (.A1(_05644_),
    .A2(_05664_),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13662_ (.A1(_05642_),
    .A2(_05665_),
    .Z(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13663_ (.A1(_05630_),
    .A2(_05666_),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13664_ (.A1(_05628_),
    .A2(_05667_),
    .Z(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13665_ (.A1(_05605_),
    .A2(_05668_),
    .Z(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13666_ (.A1(_05603_),
    .A2(_05669_),
    .Z(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13667_ (.A1(_05581_),
    .A2(_05585_),
    .A3(_05670_),
    .ZN(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13668_ (.A1(_05579_),
    .A2(_05671_),
    .ZN(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _13669_ (.A1(_05575_),
    .A2(_05576_),
    .A3(_05672_),
    .Z(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13670_ (.A1(_05575_),
    .A2(_05576_),
    .B(_05672_),
    .ZN(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13671_ (.A1(_05673_),
    .A2(_05674_),
    .Z(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13672_ (.I(\filters.low[1] ),
    .Z(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13673_ (.A1(_05676_),
    .A2(_03221_),
    .ZN(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13674_ (.A1(_03253_),
    .A2(_03378_),
    .B(_05677_),
    .ZN(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13675_ (.A1(_05675_),
    .A2(_05678_),
    .Z(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13676_ (.A1(_05574_),
    .A2(_05679_),
    .Z(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13677_ (.A1(_05573_),
    .A2(_05680_),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13678_ (.A1(_03253_),
    .A2(_05571_),
    .B(_05681_),
    .C(_03671_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13679_ (.A1(_05554_),
    .A2(_05557_),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13680_ (.A1(_05579_),
    .A2(_05671_),
    .ZN(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13681_ (.A1(_05579_),
    .A2(_05671_),
    .ZN(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13682_ (.A1(_05682_),
    .A2(_05683_),
    .B(_05684_),
    .ZN(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _13683_ (.A1(net35),
    .A2(net36),
    .B(_05558_),
    .C(_05672_),
    .ZN(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13684_ (.A1(_05594_),
    .A2(_05601_),
    .Z(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13685_ (.A1(_05591_),
    .A2(_05602_),
    .B(_05687_),
    .ZN(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13686_ (.A1(_05605_),
    .A2(_05668_),
    .ZN(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13687_ (.A1(_05603_),
    .A2(_05669_),
    .B(_05689_),
    .ZN(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13688_ (.I(_05596_),
    .Z(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13689_ (.A1(_04675_),
    .A2(_05691_),
    .A3(_05598_),
    .ZN(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13690_ (.A1(_04587_),
    .A2(_05587_),
    .A3(_05600_),
    .ZN(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13691_ (.A1(_05692_),
    .A2(_05693_),
    .Z(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13692_ (.A1(_05610_),
    .A2(_05626_),
    .ZN(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13693_ (.A1(_05608_),
    .A2(_05627_),
    .ZN(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13694_ (.A1(_05695_),
    .A2(_05696_),
    .ZN(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13695_ (.A1(_04526_),
    .A2(_05691_),
    .ZN(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13696_ (.I(_05534_),
    .Z(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13697_ (.I(_05699_),
    .Z(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13698_ (.A1(_04624_),
    .A2(_05700_),
    .A3(_05615_),
    .ZN(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13699_ (.A1(_05612_),
    .A2(_05614_),
    .B(_05701_),
    .ZN(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13700_ (.A1(_04795_),
    .A2(_05700_),
    .ZN(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13701_ (.A1(_05702_),
    .A2(_05703_),
    .ZN(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13702_ (.A1(_05698_),
    .A2(_05704_),
    .Z(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13703_ (.A1(_05697_),
    .A2(_05705_),
    .ZN(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13704_ (.A1(_05694_),
    .A2(_05706_),
    .Z(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13705_ (.I(_05628_),
    .ZN(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13706_ (.A1(_05630_),
    .A2(_05666_),
    .ZN(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13707_ (.A1(_05708_),
    .A2(_05667_),
    .B(_05709_),
    .ZN(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13708_ (.A1(_05620_),
    .A2(_05624_),
    .Z(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13709_ (.A1(_05616_),
    .A2(_05625_),
    .B(_05711_),
    .ZN(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13710_ (.I(_04474_),
    .Z(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13711_ (.A1(_04538_),
    .A2(_05713_),
    .A3(_05509_),
    .ZN(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13712_ (.A1(_05635_),
    .A2(_05714_),
    .B(_05640_),
    .ZN(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13713_ (.A1(_05633_),
    .A2(_05641_),
    .B(_05715_),
    .ZN(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13714_ (.I(_05613_),
    .Z(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13715_ (.A1(_04204_),
    .A2(_05717_),
    .ZN(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13716_ (.A1(_04325_),
    .A2(_05286_),
    .ZN(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13717_ (.I0(\filters.high[22] ),
    .I1(\filters.band[22] ),
    .S(_05207_),
    .Z(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13718_ (.A1(_04306_),
    .A2(_05720_),
    .ZN(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13719_ (.A1(_05719_),
    .A2(_05721_),
    .Z(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13720_ (.A1(_05718_),
    .A2(_05722_),
    .ZN(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13721_ (.A1(_05622_),
    .A2(_05623_),
    .Z(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13722_ (.A1(_05622_),
    .A2(_05623_),
    .Z(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13723_ (.A1(_05621_),
    .A2(_05724_),
    .B(_05725_),
    .ZN(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13724_ (.A1(_04260_),
    .A2(_05394_),
    .ZN(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13725_ (.A1(_04724_),
    .A2(_05103_),
    .ZN(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13726_ (.A1(_05540_),
    .A2(_05306_),
    .ZN(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13727_ (.A1(_05727_),
    .A2(_05728_),
    .A3(_05729_),
    .ZN(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13728_ (.A1(_05723_),
    .A2(_05726_),
    .A3(_05730_),
    .Z(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13729_ (.A1(_05716_),
    .A2(_05731_),
    .ZN(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13730_ (.A1(_05712_),
    .A2(_05732_),
    .ZN(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13731_ (.A1(_05644_),
    .A2(_05664_),
    .ZN(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13732_ (.A1(_05642_),
    .A2(_05665_),
    .B(_05734_),
    .ZN(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13733_ (.A1(_05638_),
    .A2(_05639_),
    .Z(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13734_ (.A1(_05638_),
    .A2(_05639_),
    .Z(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13735_ (.A1(_05637_),
    .A2(_05736_),
    .B(_05737_),
    .ZN(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13736_ (.A1(_05646_),
    .A2(_05647_),
    .Z(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13737_ (.A1(_05646_),
    .A2(_05647_),
    .Z(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13738_ (.A1(_05645_),
    .A2(_05739_),
    .B(_05740_),
    .ZN(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13739_ (.A1(_04398_),
    .A2(_05075_),
    .ZN(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13740_ (.A1(_04406_),
    .A2(_05496_),
    .ZN(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13741_ (.A1(_05499_),
    .A2(_05617_),
    .ZN(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13742_ (.A1(_05742_),
    .A2(_05743_),
    .A3(_05744_),
    .Z(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13743_ (.A1(_05741_),
    .A2(_05745_),
    .ZN(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13744_ (.A1(_05738_),
    .A2(_05746_),
    .ZN(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13745_ (.A1(_05658_),
    .A2(_05662_),
    .ZN(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13746_ (.A1(_05649_),
    .A2(_05663_),
    .B(_05748_),
    .ZN(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13747_ (.A1(_04474_),
    .A2(_04783_),
    .ZN(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13748_ (.I(_05491_),
    .Z(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13749_ (.A1(_03385_),
    .A2(_04372_),
    .A3(_05751_),
    .ZN(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13750_ (.A1(_03400_),
    .A2(_04431_),
    .A3(_05493_),
    .ZN(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13751_ (.A1(_05752_),
    .A2(_05753_),
    .Z(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13752_ (.A1(_05750_),
    .A2(_05754_),
    .Z(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13753_ (.A1(_05660_),
    .A2(_05661_),
    .Z(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13754_ (.A1(_05660_),
    .A2(_05661_),
    .Z(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13755_ (.A1(_05659_),
    .A2(_05756_),
    .B(_05757_),
    .ZN(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13756_ (.A1(_04322_),
    .A2(_04850_),
    .Z(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13757_ (.A1(_03335_),
    .A2(_04548_),
    .A3(_05656_),
    .ZN(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13758_ (.A1(_03352_),
    .A2(_04219_),
    .A3(_05655_),
    .ZN(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13759_ (.A1(_05760_),
    .A2(_05761_),
    .Z(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13760_ (.A1(_05759_),
    .A2(_05762_),
    .Z(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13761_ (.A1(_05758_),
    .A2(_05763_),
    .ZN(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13762_ (.A1(_05755_),
    .A2(_05764_),
    .Z(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13763_ (.A1(_05749_),
    .A2(_05765_),
    .ZN(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13764_ (.A1(_05747_),
    .A2(_05766_),
    .Z(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13765_ (.A1(_05733_),
    .A2(_05735_),
    .A3(_05767_),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13766_ (.A1(_05707_),
    .A2(_05710_),
    .A3(_05768_),
    .ZN(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13767_ (.A1(_05690_),
    .A2(_05769_),
    .Z(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13768_ (.A1(_05688_),
    .A2(_05770_),
    .Z(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13769_ (.A1(_05585_),
    .A2(_05670_),
    .ZN(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13770_ (.A1(_05585_),
    .A2(_05670_),
    .ZN(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _13771_ (.A1(_05581_),
    .A2(_05772_),
    .B(_05773_),
    .ZN(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13772_ (.A1(_05771_),
    .A2(_05774_),
    .Z(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13773_ (.A1(_05685_),
    .A2(_05686_),
    .B(_05775_),
    .ZN(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _13774_ (.A1(_05775_),
    .A2(_05685_),
    .A3(_05686_),
    .Z(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13775_ (.A1(_05776_),
    .A2(_05777_),
    .ZN(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13776_ (.I(_05778_),
    .Z(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13777_ (.I(_05779_),
    .Z(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13778_ (.A1(_03270_),
    .A2(_03377_),
    .ZN(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13779_ (.A1(_03271_),
    .A2(_03348_),
    .B(_05781_),
    .ZN(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13780_ (.I(_05782_),
    .Z(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13781_ (.A1(_05673_),
    .A2(_05674_),
    .B(_05678_),
    .ZN(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13782_ (.A1(_05673_),
    .A2(_05674_),
    .A3(_05678_),
    .ZN(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13783_ (.A1(_05564_),
    .A2(_05784_),
    .B(_05785_),
    .ZN(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13784_ (.A1(_05780_),
    .A2(_05783_),
    .A3(_05786_),
    .Z(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13785_ (.A1(_05573_),
    .A2(_05787_),
    .ZN(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13786_ (.A1(_03271_),
    .A2(_05571_),
    .B(_05788_),
    .C(_03671_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13787_ (.A1(_05697_),
    .A2(_05705_),
    .Z(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13788_ (.A1(_05694_),
    .A2(_05706_),
    .B(_05789_),
    .ZN(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13789_ (.A1(_05710_),
    .A2(_05768_),
    .Z(_05791_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13790_ (.A1(_05710_),
    .A2(_05768_),
    .Z(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13791_ (.A1(_05707_),
    .A2(_05791_),
    .B(_05792_),
    .ZN(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13792_ (.I(_05700_),
    .Z(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13793_ (.A1(_04697_),
    .A2(_05794_),
    .A3(_05702_),
    .ZN(_05795_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13794_ (.A1(_05589_),
    .A2(_05691_),
    .A3(_05704_),
    .ZN(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13795_ (.A1(_05795_),
    .A2(_05796_),
    .Z(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13796_ (.A1(_05716_),
    .A2(_05731_),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13797_ (.A1(_05712_),
    .A2(_05732_),
    .ZN(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13798_ (.A1(_05798_),
    .A2(_05799_),
    .ZN(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13799_ (.A1(_04659_),
    .A2(_05794_),
    .ZN(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13800_ (.I(_05717_),
    .Z(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13801_ (.I(_05802_),
    .Z(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13802_ (.A1(_04644_),
    .A2(_05803_),
    .A3(_05722_),
    .ZN(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13803_ (.A1(_05719_),
    .A2(_05721_),
    .B(_05804_),
    .ZN(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13804_ (.A1(_04796_),
    .A2(_05803_),
    .ZN(_05806_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13805_ (.A1(_05805_),
    .A2(_05806_),
    .ZN(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13806_ (.A1(_05801_),
    .A2(_05807_),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13807_ (.A1(_05800_),
    .A2(_05808_),
    .ZN(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13808_ (.A1(_05797_),
    .A2(_05809_),
    .Z(_05810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13809_ (.A1(_05735_),
    .A2(_05767_),
    .ZN(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13810_ (.A1(_05735_),
    .A2(_05767_),
    .ZN(_05812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13811_ (.A1(_05733_),
    .A2(_05811_),
    .B(_05812_),
    .ZN(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13812_ (.I(_05730_),
    .ZN(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13813_ (.A1(_05726_),
    .A2(_05814_),
    .ZN(_05815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13814_ (.A1(_05726_),
    .A2(_05814_),
    .ZN(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13815_ (.A1(_05723_),
    .A2(_05815_),
    .B(_05816_),
    .ZN(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13816_ (.A1(_04532_),
    .A2(_04475_),
    .A3(_05648_),
    .ZN(_05818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13817_ (.A1(_05740_),
    .A2(_05818_),
    .B(_05745_),
    .ZN(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13818_ (.A1(_05738_),
    .A2(_05746_),
    .B(_05819_),
    .ZN(_05820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13819_ (.I(_05720_),
    .Z(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13820_ (.A1(_04204_),
    .A2(_05821_),
    .ZN(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13821_ (.A1(_05211_),
    .A2(_05378_),
    .ZN(_05823_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13822_ (.I0(\filters.high[23] ),
    .I1(\filters.band[23] ),
    .S(_05207_),
    .Z(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13823_ (.A1(_04306_),
    .A2(_05824_),
    .ZN(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13824_ (.A1(_05823_),
    .A2(_05825_),
    .Z(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13825_ (.A1(_05822_),
    .A2(_05826_),
    .ZN(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _13826_ (.A1(_04271_),
    .A2(_05103_),
    .B1(_05107_),
    .B2(_04266_),
    .ZN(_05828_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13827_ (.A1(_04271_),
    .A2(_04878_),
    .A3(_04955_),
    .A4(_05107_),
    .ZN(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13828_ (.A1(_05727_),
    .A2(_05828_),
    .B(_05829_),
    .ZN(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13829_ (.A1(_04259_),
    .A2(_05286_),
    .ZN(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13830_ (.A1(_04287_),
    .A2(_05105_),
    .ZN(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13831_ (.A1(_04421_),
    .A2(_05215_),
    .ZN(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13832_ (.A1(_05831_),
    .A2(_05832_),
    .A3(_05833_),
    .ZN(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13833_ (.A1(_05830_),
    .A2(_05834_),
    .Z(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13834_ (.A1(_05827_),
    .A2(_05835_),
    .ZN(_05836_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13835_ (.A1(_05820_),
    .A2(_05836_),
    .ZN(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13836_ (.A1(_05817_),
    .A2(_05837_),
    .ZN(_05838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13837_ (.A1(_05749_),
    .A2(_05765_),
    .ZN(_05839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13838_ (.A1(_05747_),
    .A2(_05766_),
    .B(_05839_),
    .ZN(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13839_ (.A1(_05743_),
    .A2(_05744_),
    .Z(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13840_ (.A1(_05743_),
    .A2(_05744_),
    .Z(_05842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13841_ (.A1(_05742_),
    .A2(_05841_),
    .B(_05842_),
    .ZN(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13842_ (.A1(_05752_),
    .A2(_05753_),
    .Z(_05844_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13843_ (.A1(_05752_),
    .A2(_05753_),
    .Z(_05845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13844_ (.A1(_05750_),
    .A2(_05844_),
    .B(_05845_),
    .ZN(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13845_ (.A1(_04354_),
    .A2(_04955_),
    .Z(_05847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13846_ (.A1(_04480_),
    .A2(_04972_),
    .ZN(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13847_ (.A1(_04477_),
    .A2(_05076_),
    .ZN(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13848_ (.A1(_05847_),
    .A2(_05848_),
    .A3(_05849_),
    .ZN(_05850_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13849_ (.A1(_05846_),
    .A2(_05850_),
    .ZN(_05851_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13850_ (.A1(_05843_),
    .A2(_05851_),
    .ZN(_05852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13851_ (.A1(_05758_),
    .A2(_05763_),
    .ZN(_05853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13852_ (.A1(_05755_),
    .A2(_05764_),
    .B(_05853_),
    .ZN(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13853_ (.A1(_04473_),
    .A2(_04788_),
    .ZN(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13854_ (.A1(_04531_),
    .A2(_05751_),
    .ZN(_05856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13855_ (.I(_05493_),
    .Z(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13856_ (.A1(_04783_),
    .A2(_05857_),
    .ZN(_05858_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13857_ (.A1(_05855_),
    .A2(_05856_),
    .A3(_05858_),
    .Z(_05859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13858_ (.A1(_05760_),
    .A2(_05761_),
    .ZN(_05860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13859_ (.A1(_05759_),
    .A2(_05762_),
    .B(_05860_),
    .ZN(_05861_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13860_ (.A1(_04427_),
    .A2(_04850_),
    .Z(_05862_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13861_ (.A1(_03351_),
    .A2(_04218_),
    .A3(_05651_),
    .ZN(_05863_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13862_ (.A1(_03366_),
    .A2(_04885_),
    .A3(_05654_),
    .ZN(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13863_ (.A1(_05863_),
    .A2(_05864_),
    .Z(_05865_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13864_ (.A1(_05862_),
    .A2(_05865_),
    .ZN(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13865_ (.A1(_05861_),
    .A2(_05866_),
    .ZN(_05867_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13866_ (.A1(_05859_),
    .A2(_05867_),
    .Z(_05868_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13867_ (.A1(_05854_),
    .A2(_05868_),
    .ZN(_05869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13868_ (.A1(_05852_),
    .A2(_05869_),
    .Z(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13869_ (.A1(_05838_),
    .A2(_05840_),
    .A3(_05870_),
    .ZN(_05871_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13870_ (.A1(_05810_),
    .A2(_05813_),
    .A3(_05871_),
    .ZN(_05872_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _13871_ (.A1(_05790_),
    .A2(_05793_),
    .A3(_05872_),
    .ZN(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13872_ (.A1(_05690_),
    .A2(_05769_),
    .ZN(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13873_ (.A1(_05688_),
    .A2(_05770_),
    .B(_05874_),
    .ZN(_05875_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13874_ (.A1(_05873_),
    .A2(_05875_),
    .Z(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13875_ (.A1(_05771_),
    .A2(_05774_),
    .ZN(_05877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _13876_ (.A1(_05776_),
    .A2(_05877_),
    .ZN(_05878_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _13877_ (.A1(_05878_),
    .A2(_05876_),
    .ZN(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13878_ (.I(_03378_),
    .Z(_05880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13879_ (.A1(_03284_),
    .A2(_03222_),
    .ZN(_05881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13880_ (.A1(_03286_),
    .A2(_05880_),
    .B(_05881_),
    .ZN(_05882_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13881_ (.A1(_05879_),
    .A2(_05882_),
    .Z(_05883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13882_ (.A1(_05780_),
    .A2(_05783_),
    .ZN(_05884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13883_ (.A1(_05574_),
    .A2(_05679_),
    .ZN(_05885_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13884_ (.A1(_05785_),
    .A2(_05885_),
    .Z(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13885_ (.A1(_05780_),
    .A2(_05783_),
    .ZN(_05887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13886_ (.A1(_05884_),
    .A2(_05886_),
    .B(_05887_),
    .ZN(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13887_ (.A1(_05883_),
    .A2(_05888_),
    .Z(_05889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13888_ (.A1(_05573_),
    .A2(_05889_),
    .ZN(_05890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13889_ (.A1(_03286_),
    .A2(_05571_),
    .B(_05890_),
    .C(_03671_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13890_ (.A1(_05879_),
    .A2(_05882_),
    .ZN(_05891_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13891_ (.A1(_05778_),
    .A2(_05783_),
    .Z(_05892_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13892_ (.A1(_05778_),
    .A2(_05782_),
    .Z(_05893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13893_ (.A1(_05892_),
    .A2(_05786_),
    .B(_05893_),
    .ZN(_05894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13894_ (.A1(_05882_),
    .A2(_05879_),
    .ZN(_05895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13895_ (.A1(_05891_),
    .A2(_05894_),
    .B(_05895_),
    .ZN(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13896_ (.A1(_05558_),
    .A2(_05672_),
    .ZN(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13897_ (.A1(_05775_),
    .A2(_05897_),
    .A3(_05876_),
    .ZN(_05898_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _13898_ (.A1(_05775_),
    .A2(_05685_),
    .A3(_05876_),
    .ZN(_05899_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13899_ (.A1(_05771_),
    .A2(_05774_),
    .Z(_05900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13900_ (.A1(_05873_),
    .A2(_05875_),
    .ZN(_05901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13901_ (.A1(_05873_),
    .A2(_05875_),
    .ZN(_05902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13902_ (.A1(_05900_),
    .A2(_05901_),
    .B(_05902_),
    .ZN(_05903_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _13903_ (.A1(_05461_),
    .A2(_05898_),
    .B(_05899_),
    .C(_05903_),
    .ZN(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13904_ (.A1(_05800_),
    .A2(_05808_),
    .Z(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13905_ (.A1(_05797_),
    .A2(_05809_),
    .B(_05905_),
    .ZN(_05906_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13906_ (.A1(_05813_),
    .A2(_05871_),
    .Z(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13907_ (.A1(_05813_),
    .A2(_05871_),
    .Z(_05908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13908_ (.A1(_05810_),
    .A2(_05907_),
    .B(_05908_),
    .ZN(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13909_ (.I(_05803_),
    .Z(_05910_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13910_ (.A1(_04675_),
    .A2(_05910_),
    .A3(_05805_),
    .ZN(_05911_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13911_ (.A1(_04660_),
    .A2(_05794_),
    .A3(_05807_),
    .ZN(_05912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13912_ (.A1(_05911_),
    .A2(_05912_),
    .Z(_05913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13913_ (.A1(_05820_),
    .A2(_05836_),
    .ZN(_05914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13914_ (.A1(_05817_),
    .A2(_05837_),
    .ZN(_05915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13915_ (.A1(_05914_),
    .A2(_05915_),
    .ZN(_05916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13916_ (.A1(_04658_),
    .A2(_05910_),
    .ZN(_05917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13917_ (.I(_05821_),
    .Z(_05918_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13918_ (.A1(_04606_),
    .A2(_05918_),
    .A3(_05826_),
    .ZN(_05919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13919_ (.A1(_05823_),
    .A2(_05825_),
    .B(_05919_),
    .ZN(_05920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13920_ (.I(_05918_),
    .Z(_05921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13921_ (.A1(_04795_),
    .A2(_05921_),
    .ZN(_05922_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13922_ (.A1(_05920_),
    .A2(_05922_),
    .ZN(_05923_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13923_ (.A1(_05917_),
    .A2(_05923_),
    .Z(_05924_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13924_ (.A1(_05916_),
    .A2(_05924_),
    .ZN(_05925_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13925_ (.A1(_05913_),
    .A2(_05925_),
    .Z(_05926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13926_ (.A1(_05840_),
    .A2(_05870_),
    .ZN(_05927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13927_ (.A1(_05840_),
    .A2(_05870_),
    .ZN(_05928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13928_ (.A1(_05838_),
    .A2(_05927_),
    .B(_05928_),
    .ZN(_05929_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13929_ (.A1(_05830_),
    .A2(_05834_),
    .Z(_05930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13930_ (.A1(_05827_),
    .A2(_05835_),
    .B(_05930_),
    .ZN(_05931_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13931_ (.A1(_05713_),
    .A2(_04799_),
    .A3(_05754_),
    .ZN(_05932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13932_ (.A1(_05845_),
    .A2(_05932_),
    .B(_05850_),
    .ZN(_05933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13933_ (.A1(_05843_),
    .A2(_05851_),
    .B(_05933_),
    .ZN(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13934_ (.A1(_04551_),
    .A2(_05824_),
    .ZN(_05935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13935_ (.A1(_04227_),
    .A2(_05533_),
    .ZN(_05936_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13936_ (.I0(\filters.high[24] ),
    .I1(\filters.band[24] ),
    .S(_03190_),
    .Z(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13937_ (.A1(_04513_),
    .A2(_05937_),
    .ZN(_05938_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13938_ (.A1(_05936_),
    .A2(_05938_),
    .Z(_05939_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13939_ (.A1(_05935_),
    .A2(_05939_),
    .ZN(_05940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13940_ (.I(_04250_),
    .Z(_05941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13941_ (.A1(_04724_),
    .A2(_05305_),
    .B1(_05395_),
    .B2(_05941_),
    .ZN(_05942_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13942_ (.A1(_04724_),
    .A2(_05941_),
    .A3(_05305_),
    .A4(_05216_),
    .ZN(_05943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13943_ (.A1(_05831_),
    .A2(_05942_),
    .B(_05943_),
    .ZN(_05944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13944_ (.A1(_04734_),
    .A2(_05529_),
    .ZN(_05945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13945_ (.A1(_04270_),
    .A2(_05215_),
    .ZN(_05946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13946_ (.I(_05286_),
    .Z(_05947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13947_ (.A1(_04878_),
    .A2(_05947_),
    .ZN(_05948_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13948_ (.A1(_05945_),
    .A2(_05946_),
    .A3(_05948_),
    .ZN(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13949_ (.A1(_05944_),
    .A2(_05949_),
    .Z(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13950_ (.A1(_05940_),
    .A2(_05950_),
    .ZN(_05951_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13951_ (.A1(_05934_),
    .A2(_05951_),
    .ZN(_05952_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13952_ (.A1(_05931_),
    .A2(_05952_),
    .ZN(_05953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13953_ (.A1(_05854_),
    .A2(_05868_),
    .ZN(_05954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13954_ (.A1(_05852_),
    .A2(_05869_),
    .B(_05954_),
    .ZN(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13955_ (.A1(_05848_),
    .A2(_05849_),
    .ZN(_05956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13956_ (.A1(_05848_),
    .A2(_05849_),
    .ZN(_05957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13957_ (.A1(_05847_),
    .A2(_05956_),
    .B(_05957_),
    .ZN(_05958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13958_ (.I(_05491_),
    .Z(_05959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13959_ (.A1(_04531_),
    .A2(_05959_),
    .B1(_04837_),
    .B2(_04783_),
    .ZN(_05960_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _13960_ (.A1(_04531_),
    .A2(_04798_),
    .A3(_05751_),
    .A4(_04837_),
    .ZN(_05961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13961_ (.A1(_05855_),
    .A2(_05960_),
    .B(_05961_),
    .ZN(_05962_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13962_ (.A1(_04398_),
    .A2(_05106_),
    .Z(_05963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13963_ (.A1(_04406_),
    .A2(_05075_),
    .ZN(_05964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13964_ (.A1(_04346_),
    .A2(_05103_),
    .ZN(_05965_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13965_ (.A1(_05963_),
    .A2(_05964_),
    .A3(_05965_),
    .Z(_05966_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13966_ (.A1(_05962_),
    .A2(_05966_),
    .ZN(_05967_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13967_ (.A1(_05958_),
    .A2(_05967_),
    .ZN(_05968_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13968_ (.A1(_05861_),
    .A2(_05866_),
    .Z(_05969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13969_ (.A1(_05859_),
    .A2(_05867_),
    .B(_05969_),
    .ZN(_05970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13970_ (.A1(_05863_),
    .A2(_05864_),
    .ZN(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13971_ (.A1(_05862_),
    .A2(_05865_),
    .B(_05971_),
    .ZN(_05972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13972_ (.A1(_04303_),
    .A2(_05651_),
    .ZN(_05973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13973_ (.A1(_04426_),
    .A2(_05654_),
    .ZN(_05974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13974_ (.A1(_04433_),
    .A2(_04849_),
    .ZN(_05975_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13975_ (.A1(_05973_),
    .A2(_05974_),
    .A3(_05975_),
    .Z(_05976_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13976_ (.A1(_05972_),
    .A2(_05976_),
    .ZN(_05977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13977_ (.A1(_04472_),
    .A2(_05617_),
    .ZN(_05978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13978_ (.A1(_04782_),
    .A2(_05491_),
    .ZN(_05979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13979_ (.A1(_04788_),
    .A2(_05493_),
    .ZN(_05980_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _13980_ (.A1(_05978_),
    .A2(_05979_),
    .A3(_05980_),
    .Z(_05981_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13981_ (.A1(_05977_),
    .A2(_05981_),
    .Z(_05982_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13982_ (.A1(_05970_),
    .A2(_05982_),
    .ZN(_05983_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13983_ (.A1(_05968_),
    .A2(_05983_),
    .Z(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13984_ (.A1(_05953_),
    .A2(_05955_),
    .A3(_05984_),
    .ZN(_05985_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _13985_ (.A1(_05926_),
    .A2(_05929_),
    .A3(_05985_),
    .ZN(_05986_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13986_ (.A1(_05909_),
    .A2(_05986_),
    .Z(_05987_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _13987_ (.A1(_05906_),
    .A2(_05987_),
    .ZN(_05988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13988_ (.A1(_05793_),
    .A2(_05872_),
    .ZN(_05989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13989_ (.A1(_05793_),
    .A2(_05872_),
    .ZN(_05990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _13990_ (.A1(_05790_),
    .A2(_05989_),
    .B(_05990_),
    .ZN(_05991_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13991_ (.A1(_05988_),
    .A2(_05991_),
    .Z(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _13992_ (.A1(_05904_),
    .A2(_05992_),
    .Z(_05993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13993_ (.I(\filters.low[4] ),
    .Z(_05994_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13994_ (.A1(_05994_),
    .A2(_03473_),
    .ZN(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13995_ (.A1(_03301_),
    .A2(_03473_),
    .B(_05995_),
    .ZN(_05996_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13996_ (.A1(_05993_),
    .A2(_05996_),
    .Z(_05997_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13997_ (.A1(_05896_),
    .A2(_05997_),
    .Z(_05998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13998_ (.A1(\filters.band[4] ),
    .A2(_05567_),
    .B(_03753_),
    .ZN(_05999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13999_ (.A1(_04189_),
    .A2(_05998_),
    .B(_05999_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14000_ (.I(_05569_),
    .Z(_06000_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14001_ (.A1(_05916_),
    .A2(_05924_),
    .Z(_06001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14002_ (.A1(_05913_),
    .A2(_05925_),
    .B(_06001_),
    .ZN(_06002_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14003_ (.A1(_05929_),
    .A2(_05985_),
    .Z(_06003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14004_ (.A1(_05929_),
    .A2(_05985_),
    .Z(_06004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14005_ (.A1(_05926_),
    .A2(_06003_),
    .B(_06004_),
    .ZN(_06005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14006_ (.I(_05921_),
    .Z(_06006_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14007_ (.A1(_05586_),
    .A2(_06006_),
    .A3(_05920_),
    .ZN(_06007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14008_ (.I(_04660_),
    .Z(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14009_ (.A1(_06008_),
    .A2(_05910_),
    .A3(_05923_),
    .ZN(_06009_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14010_ (.A1(_06007_),
    .A2(_06009_),
    .Z(_06010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14011_ (.A1(_05934_),
    .A2(_05951_),
    .ZN(_06011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14012_ (.A1(_05931_),
    .A2(_05952_),
    .ZN(_06012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14013_ (.A1(_06011_),
    .A2(_06012_),
    .ZN(_06013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14014_ (.A1(_04659_),
    .A2(_05921_),
    .ZN(_06014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14015_ (.I(_05824_),
    .Z(_06015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14016_ (.I(_06015_),
    .Z(_06016_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14017_ (.A1(_04644_),
    .A2(_06016_),
    .A3(_05939_),
    .ZN(_06017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14018_ (.A1(_05936_),
    .A2(_05938_),
    .B(_06017_),
    .ZN(_06018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14019_ (.A1(_04524_),
    .A2(_06016_),
    .ZN(_06019_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14020_ (.A1(_06018_),
    .A2(_06019_),
    .ZN(_06020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14021_ (.A1(_06014_),
    .A2(_06020_),
    .Z(_06021_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14022_ (.A1(_06013_),
    .A2(_06021_),
    .ZN(_06022_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14023_ (.A1(_06010_),
    .A2(_06022_),
    .Z(_06023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14024_ (.A1(_05955_),
    .A2(_05984_),
    .ZN(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14025_ (.A1(_05955_),
    .A2(_05984_),
    .ZN(_06025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14026_ (.A1(_05953_),
    .A2(_06024_),
    .B(_06025_),
    .ZN(_06026_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14027_ (.A1(_05944_),
    .A2(_05949_),
    .Z(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14028_ (.A1(_05940_),
    .A2(_05950_),
    .B(_06027_),
    .ZN(_06028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14029_ (.A1(_05962_),
    .A2(_05966_),
    .ZN(_06029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14030_ (.A1(_05958_),
    .A2(_05967_),
    .B(_06029_),
    .ZN(_06030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14031_ (.I(_05937_),
    .Z(_06031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14032_ (.A1(_04555_),
    .A2(_06031_),
    .ZN(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14033_ (.A1(_05211_),
    .A2(_05613_),
    .ZN(_06033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14034_ (.I0(\filters.high[25] ),
    .I1(\filters.band[25] ),
    .S(_03190_),
    .Z(_06034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14035_ (.A1(_04214_),
    .A2(_06034_),
    .ZN(_06035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14036_ (.A1(_06033_),
    .A2(_06035_),
    .Z(_06036_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14037_ (.A1(_06032_),
    .A2(_06036_),
    .ZN(_06037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14038_ (.A1(_05538_),
    .A2(_05395_),
    .B1(_05474_),
    .B2(_05941_),
    .ZN(_06038_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _14039_ (.A1(_05538_),
    .A2(_05941_),
    .A3(_05216_),
    .A4(_05947_),
    .ZN(_06039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14040_ (.A1(_05945_),
    .A2(_06038_),
    .B(_06039_),
    .ZN(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _14041_ (.A1(_04759_),
    .A2(_05374_),
    .ZN(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14042_ (.A1(_04506_),
    .A2(_05378_),
    .ZN(_06042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14043_ (.A1(_04260_),
    .A2(_05533_),
    .ZN(_06043_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14044_ (.A1(_06041_),
    .A2(_06042_),
    .A3(_06043_),
    .ZN(_06044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14045_ (.A1(_06040_),
    .A2(_06044_),
    .Z(_06045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14046_ (.A1(_06037_),
    .A2(_06045_),
    .Z(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14047_ (.A1(_06030_),
    .A2(_06046_),
    .ZN(_06047_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14048_ (.A1(_06028_),
    .A2(_06047_),
    .ZN(_06048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14049_ (.A1(_05970_),
    .A2(_05982_),
    .ZN(_06049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14050_ (.A1(_05968_),
    .A2(_05983_),
    .B(_06049_),
    .ZN(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14051_ (.A1(_05972_),
    .A2(_05976_),
    .Z(_06051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14052_ (.A1(_05977_),
    .A2(_05981_),
    .B(_06051_),
    .ZN(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14053_ (.A1(_04427_),
    .A2(_05655_),
    .B1(_05656_),
    .B2(_04303_),
    .ZN(_06053_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _14054_ (.A1(_04304_),
    .A2(_04427_),
    .A3(_05655_),
    .A4(_05656_),
    .ZN(_06054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14055_ (.A1(_06053_),
    .A2(_05975_),
    .B(_06054_),
    .ZN(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14056_ (.A1(_03384_),
    .A2(_04371_),
    .A3(_05135_),
    .ZN(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14057_ (.A1(net54),
    .A2(_04431_),
    .A3(_04911_),
    .ZN(_06057_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14058_ (.A1(_06056_),
    .A2(_06057_),
    .ZN(_06058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14059_ (.A1(_04780_),
    .A2(_04914_),
    .ZN(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14060_ (.A1(_06058_),
    .A2(_06059_),
    .Z(_06060_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14061_ (.A1(_06055_),
    .A2(_06060_),
    .ZN(_06061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14062_ (.A1(_04824_),
    .A2(_04893_),
    .ZN(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14063_ (.A1(_05496_),
    .A2(_04856_),
    .ZN(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14064_ (.A1(_05212_),
    .A2(_05256_),
    .ZN(_06064_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14065_ (.A1(_06062_),
    .A2(_06063_),
    .A3(_06064_),
    .Z(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14066_ (.A1(_06061_),
    .A2(_06065_),
    .Z(_06066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14067_ (.A1(_06052_),
    .A2(_06066_),
    .Z(_06067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14068_ (.A1(_05964_),
    .A2(_05965_),
    .ZN(_06068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14069_ (.A1(_05964_),
    .A2(_05965_),
    .ZN(_06069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14070_ (.A1(_05963_),
    .A2(_06068_),
    .B(_06069_),
    .ZN(_06070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14071_ (.A1(_04798_),
    .A2(_05492_),
    .B1(_04836_),
    .B2(_05539_),
    .ZN(_06071_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _14072_ (.A1(_04782_),
    .A2(_05539_),
    .A3(_05492_),
    .A4(_04836_),
    .ZN(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14073_ (.A1(_05978_),
    .A2(_06071_),
    .B(_06072_),
    .ZN(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14074_ (.A1(_04479_),
    .A2(_05102_),
    .ZN(_06074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14075_ (.A1(_04752_),
    .A2(_05106_),
    .ZN(_06075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14076_ (.A1(_04354_),
    .A2(_05394_),
    .ZN(_06076_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14077_ (.A1(_06074_),
    .A2(_06075_),
    .A3(_06076_),
    .Z(_06077_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14078_ (.A1(_06073_),
    .A2(_06077_),
    .Z(_06078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14079_ (.A1(_06070_),
    .A2(_06078_),
    .Z(_06079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14080_ (.A1(_06067_),
    .A2(_06079_),
    .Z(_06080_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14081_ (.A1(_06050_),
    .A2(_06080_),
    .ZN(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14082_ (.A1(_06048_),
    .A2(_06081_),
    .Z(_06082_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14083_ (.A1(_06023_),
    .A2(_06026_),
    .A3(_06082_),
    .ZN(_06083_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14084_ (.A1(_06002_),
    .A2(_06005_),
    .A3(_06083_),
    .ZN(_06084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14085_ (.A1(_05909_),
    .A2(_05986_),
    .ZN(_06085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14086_ (.A1(_05906_),
    .A2(_05987_),
    .B(_06085_),
    .ZN(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14087_ (.A1(_06084_),
    .A2(_06086_),
    .Z(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _14088_ (.A1(_05988_),
    .A2(_05991_),
    .ZN(_06088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14089_ (.A1(_05904_),
    .A2(_05992_),
    .B(_06088_),
    .ZN(_06089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14090_ (.A1(_06087_),
    .A2(_06089_),
    .Z(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14091_ (.I(_03377_),
    .Z(_06091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14092_ (.I(_06091_),
    .Z(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14093_ (.A1(_03312_),
    .A2(_03379_),
    .ZN(_06093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14094_ (.A1(_03316_),
    .A2(_06092_),
    .B(_06093_),
    .ZN(_06094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14095_ (.A1(_06090_),
    .A2(_06094_),
    .ZN(_06095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14096_ (.A1(_06090_),
    .A2(_06094_),
    .Z(_06096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14097_ (.A1(_06095_),
    .A2(_06096_),
    .ZN(_06097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _14098_ (.I(_03474_),
    .Z(_06098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _14099_ (.A1(_03301_),
    .A2(_06098_),
    .B(_05993_),
    .C(_05995_),
    .ZN(_06099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14100_ (.A1(_05883_),
    .A2(_05888_),
    .ZN(_06100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14101_ (.A1(_05895_),
    .A2(_06100_),
    .B(_05997_),
    .ZN(_06101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14102_ (.A1(_06099_),
    .A2(_06101_),
    .ZN(_06102_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14103_ (.A1(_06097_),
    .A2(_06102_),
    .ZN(_06103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14104_ (.A1(_06000_),
    .A2(_06103_),
    .ZN(_06104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14105_ (.I(_01827_),
    .Z(_06105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14106_ (.A1(_03316_),
    .A2(_05571_),
    .B(_06104_),
    .C(_06105_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14107_ (.I(_05570_),
    .Z(_06106_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14108_ (.A1(_06013_),
    .A2(_06021_),
    .Z(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14109_ (.A1(_06010_),
    .A2(_06022_),
    .B(_06107_),
    .ZN(_06108_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14110_ (.A1(_06026_),
    .A2(_06082_),
    .Z(_06109_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14111_ (.A1(_06026_),
    .A2(_06082_),
    .Z(_06110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14112_ (.A1(_06023_),
    .A2(_06109_),
    .B(_06110_),
    .ZN(_06111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14113_ (.I(_06016_),
    .Z(_06112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14114_ (.A1(_04697_),
    .A2(_06112_),
    .A3(_06018_),
    .ZN(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14115_ (.A1(_04669_),
    .A2(_06006_),
    .A3(_06020_),
    .ZN(_06114_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14116_ (.A1(_06113_),
    .A2(_06114_),
    .Z(_06115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14117_ (.A1(_06028_),
    .A2(_06047_),
    .ZN(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14118_ (.A1(_06030_),
    .A2(_06046_),
    .B(_06116_),
    .ZN(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14119_ (.A1(_04586_),
    .A2(_06112_),
    .ZN(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14120_ (.I(_06031_),
    .Z(_06119_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14121_ (.A1(_04625_),
    .A2(_06119_),
    .A3(_06036_),
    .ZN(_06120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14122_ (.A1(_06033_),
    .A2(_06035_),
    .B(_06120_),
    .ZN(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14123_ (.A1(_04672_),
    .A2(_06119_),
    .ZN(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14124_ (.A1(_06121_),
    .A2(_06122_),
    .ZN(_06123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14125_ (.A1(_06118_),
    .A2(_06123_),
    .Z(_06124_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14126_ (.A1(_06117_),
    .A2(_06124_),
    .ZN(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14127_ (.A1(_06115_),
    .A2(_06125_),
    .Z(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14128_ (.A1(_06050_),
    .A2(_06080_),
    .ZN(_06127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14129_ (.A1(_06048_),
    .A2(_06081_),
    .B(_06127_),
    .ZN(_06128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14130_ (.A1(_06052_),
    .A2(_06066_),
    .Z(_06129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14131_ (.A1(_06067_),
    .A2(_06079_),
    .B(_06129_),
    .ZN(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14132_ (.A1(_06055_),
    .A2(_06060_),
    .ZN(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14133_ (.A1(_06061_),
    .A2(_06065_),
    .B(_06131_),
    .ZN(_06132_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14134_ (.A1(_06056_),
    .A2(_06057_),
    .Z(_06133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14135_ (.A1(_06058_),
    .A2(_06059_),
    .B(_06133_),
    .ZN(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _14136_ (.A1(net55),
    .A2(_04430_),
    .A3(_05134_),
    .ZN(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _14137_ (.A1(_03415_),
    .A2(_04514_),
    .A3(_04910_),
    .ZN(_06136_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14138_ (.A1(_06135_),
    .A2(_06136_),
    .ZN(_06137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14139_ (.A1(_04740_),
    .A2(_04848_),
    .ZN(_06138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14140_ (.A1(_06137_),
    .A2(_06138_),
    .ZN(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14141_ (.A1(_06134_),
    .A2(_06139_),
    .ZN(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14142_ (.A1(_04771_),
    .A2(_04814_),
    .ZN(_06141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14143_ (.A1(_04834_),
    .A2(_04892_),
    .ZN(_06142_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14144_ (.A1(_06141_),
    .A2(_06142_),
    .ZN(_06143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _14145_ (.A1(_04472_),
    .A2(_04955_),
    .ZN(_06144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14146_ (.A1(_06143_),
    .A2(_06144_),
    .Z(_06145_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14147_ (.A1(_06140_),
    .A2(_06145_),
    .Z(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14148_ (.A1(_06132_),
    .A2(_06146_),
    .Z(_06147_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14149_ (.A1(_06074_),
    .A2(_06075_),
    .Z(_06148_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14150_ (.A1(_06074_),
    .A2(_06075_),
    .Z(_06149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14151_ (.A1(_06148_),
    .A2(_06076_),
    .B(_06149_),
    .ZN(_06150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14152_ (.A1(_06063_),
    .A2(_06064_),
    .Z(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14153_ (.A1(_06063_),
    .A2(_06064_),
    .Z(_06152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14154_ (.A1(_06062_),
    .A2(_06151_),
    .B(_06152_),
    .ZN(_06153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14155_ (.A1(_04405_),
    .A2(_05105_),
    .ZN(_06154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14156_ (.A1(_04344_),
    .A2(_05214_),
    .ZN(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14157_ (.A1(_05150_),
    .A2(_05374_),
    .ZN(_06156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14158_ (.A1(_06154_),
    .A2(_06155_),
    .A3(_06156_),
    .ZN(_06157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14159_ (.A1(_06153_),
    .A2(_06157_),
    .Z(_06158_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14160_ (.A1(_06150_),
    .A2(_06158_),
    .Z(_06159_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14161_ (.A1(_06147_),
    .A2(_06159_),
    .ZN(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14162_ (.A1(_06130_),
    .A2(_06160_),
    .ZN(_06161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14163_ (.A1(_06040_),
    .A2(_06044_),
    .ZN(_06162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14164_ (.A1(_06037_),
    .A2(_06045_),
    .ZN(_06163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14165_ (.A1(_06162_),
    .A2(_06163_),
    .ZN(_06164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14166_ (.I(_06077_),
    .ZN(_06165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14167_ (.A1(_06070_),
    .A2(_06078_),
    .ZN(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14168_ (.A1(_06073_),
    .A2(_06165_),
    .B(_06166_),
    .ZN(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14169_ (.A1(_04555_),
    .A2(_06034_),
    .ZN(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14170_ (.A1(_05211_),
    .A2(_05720_),
    .ZN(_06169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14171_ (.A1(\filters.band[26] ),
    .A2(_04214_),
    .ZN(_06170_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14172_ (.A1(_06169_),
    .A2(_06170_),
    .Z(_06171_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14173_ (.A1(_06168_),
    .A2(_06171_),
    .ZN(_06172_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14174_ (.A1(_06041_),
    .A2(_06042_),
    .Z(_06173_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14175_ (.A1(_06041_),
    .A2(_06042_),
    .Z(_06174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14176_ (.A1(_06173_),
    .A2(_06043_),
    .B(_06174_),
    .ZN(_06175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14177_ (.A1(_05097_),
    .A2(_05377_),
    .ZN(_06176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14178_ (.A1(_04264_),
    .A2(_05533_),
    .ZN(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14179_ (.A1(_06176_),
    .A2(_06177_),
    .Z(_06178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14180_ (.A1(_04260_),
    .A2(_05613_),
    .ZN(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14181_ (.A1(_06178_),
    .A2(_06179_),
    .ZN(_06180_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14182_ (.A1(_06175_),
    .A2(_06180_),
    .Z(_06181_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14183_ (.A1(_06172_),
    .A2(_06181_),
    .ZN(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14184_ (.A1(_06167_),
    .A2(_06182_),
    .Z(_06183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14185_ (.A1(_06164_),
    .A2(_06183_),
    .ZN(_06184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14186_ (.A1(_06161_),
    .A2(_06184_),
    .Z(_06185_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14187_ (.A1(_06128_),
    .A2(_06185_),
    .Z(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14188_ (.A1(_06126_),
    .A2(_06186_),
    .ZN(_06187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14189_ (.A1(_06111_),
    .A2(_06187_),
    .Z(_06188_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14190_ (.A1(_06108_),
    .A2(_06188_),
    .ZN(_06189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14191_ (.A1(_06005_),
    .A2(_06083_),
    .ZN(_06190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14192_ (.A1(_06005_),
    .A2(_06083_),
    .ZN(_06191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14193_ (.A1(_06002_),
    .A2(_06190_),
    .B(_06191_),
    .ZN(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _14194_ (.A1(_06189_),
    .A2(_06192_),
    .Z(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14195_ (.A1(_05992_),
    .A2(_06087_),
    .ZN(_06194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14196_ (.I(_06194_),
    .ZN(_06195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14197_ (.A1(_06084_),
    .A2(_06086_),
    .ZN(_06196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14198_ (.A1(_06084_),
    .A2(_06086_),
    .ZN(_06197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14199_ (.A1(_06088_),
    .A2(_06196_),
    .B(_06197_),
    .ZN(_06198_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14200_ (.I(_06198_),
    .ZN(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14201_ (.A1(_05904_),
    .A2(_06195_),
    .B(_06199_),
    .ZN(_06200_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14202_ (.A1(_06193_),
    .A2(_06200_),
    .Z(_06201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _14203_ (.I(_06091_),
    .Z(_06202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14204_ (.A1(_03331_),
    .A2(_05880_),
    .ZN(_06203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _14205_ (.A1(_03332_),
    .A2(_06202_),
    .B(_06203_),
    .ZN(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14206_ (.A1(_06201_),
    .A2(_06204_),
    .Z(_06205_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _14207_ (.I(_06095_),
    .ZN(_06206_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _14208_ (.A1(_05997_),
    .A2(_06095_),
    .A3(_06096_),
    .ZN(_06207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _14209_ (.A1(_06099_),
    .A2(_06206_),
    .B1(_06207_),
    .B2(_05896_),
    .C(_06096_),
    .ZN(_06208_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14210_ (.A1(_06205_),
    .A2(_06208_),
    .ZN(_06209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14211_ (.A1(_06000_),
    .A2(_06209_),
    .ZN(_06210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14212_ (.A1(_03332_),
    .A2(_06106_),
    .B(_06210_),
    .C(_06105_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14213_ (.A1(_06117_),
    .A2(_06124_),
    .Z(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14214_ (.A1(_06115_),
    .A2(_06125_),
    .B(_06211_),
    .ZN(_06212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14215_ (.A1(_06128_),
    .A2(_06185_),
    .ZN(_06213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14216_ (.A1(_06126_),
    .A2(_06186_),
    .ZN(_06214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14217_ (.A1(_06213_),
    .A2(_06214_),
    .ZN(_06215_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14218_ (.A1(_06130_),
    .A2(_06160_),
    .Z(_06216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14219_ (.A1(_06161_),
    .A2(_06184_),
    .B(_06216_),
    .ZN(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14220_ (.A1(_06132_),
    .A2(_06146_),
    .ZN(_06218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14221_ (.A1(_06147_),
    .A2(_06159_),
    .ZN(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _14222_ (.A1(_06218_),
    .A2(_06219_),
    .ZN(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14223_ (.I(_06139_),
    .ZN(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14224_ (.A1(_06134_),
    .A2(_06221_),
    .ZN(_06222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14225_ (.A1(_06140_),
    .A2(_06145_),
    .ZN(_06223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14226_ (.A1(_06222_),
    .A2(_06223_),
    .ZN(_06224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14227_ (.A1(_06135_),
    .A2(_06136_),
    .ZN(_06225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14228_ (.A1(_06137_),
    .A2(_06138_),
    .ZN(_06226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14229_ (.A1(_06225_),
    .A2(_06226_),
    .ZN(_06227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14230_ (.A1(_04780_),
    .A2(_05514_),
    .ZN(_06228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14231_ (.A1(_04768_),
    .A2(_05654_),
    .ZN(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14232_ (.A1(_06228_),
    .A2(_06229_),
    .ZN(_06230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14233_ (.A1(_04972_),
    .A2(_04849_),
    .ZN(_06231_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14234_ (.A1(_06230_),
    .A2(_06231_),
    .ZN(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14235_ (.A1(_06227_),
    .A2(_06232_),
    .ZN(_06233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14236_ (.A1(_05492_),
    .A2(_05076_),
    .ZN(_06234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14237_ (.A1(_04836_),
    .A2(_05119_),
    .ZN(_06235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14238_ (.A1(_04925_),
    .A2(_05209_),
    .ZN(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14239_ (.A1(_06234_),
    .A2(_06235_),
    .A3(_06236_),
    .ZN(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14240_ (.A1(_06233_),
    .A2(_06237_),
    .Z(_06238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14241_ (.A1(_06224_),
    .A2(_06238_),
    .Z(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14242_ (.A1(_06154_),
    .A2(_06155_),
    .Z(_06240_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14243_ (.A1(_06154_),
    .A2(_06155_),
    .Z(_06241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14244_ (.A1(_06240_),
    .A2(_06156_),
    .B(_06241_),
    .ZN(_06242_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14245_ (.A1(_06141_),
    .A2(_06142_),
    .Z(_06243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14246_ (.A1(_06143_),
    .A2(_06144_),
    .B(_06243_),
    .ZN(_06244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14247_ (.A1(_04354_),
    .A2(_05530_),
    .ZN(_06245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14248_ (.A1(_04480_),
    .A2(_05394_),
    .ZN(_06246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14249_ (.A1(_05499_),
    .A2(_05947_),
    .ZN(_06247_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14250_ (.A1(_06246_),
    .A2(_06247_),
    .Z(_06248_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14251_ (.A1(_06245_),
    .A2(_06248_),
    .ZN(_06249_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14252_ (.A1(_06244_),
    .A2(_06249_),
    .Z(_06250_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14253_ (.A1(_06242_),
    .A2(_06250_),
    .Z(_06251_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14254_ (.A1(_06239_),
    .A2(_06251_),
    .Z(_06252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14255_ (.A1(_06220_),
    .A2(_06252_),
    .Z(_06253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14256_ (.A1(_06175_),
    .A2(_06180_),
    .ZN(_06254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14257_ (.A1(_06172_),
    .A2(_06181_),
    .ZN(_06255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14258_ (.A1(_06254_),
    .A2(_06255_),
    .ZN(_06256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14259_ (.A1(_06153_),
    .A2(_06157_),
    .ZN(_06257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14260_ (.A1(_06150_),
    .A2(_06158_),
    .ZN(_06258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _14261_ (.A1(_06257_),
    .A2(_06258_),
    .ZN(_06259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14262_ (.A1(\filters.band[26] ),
    .A2(_04624_),
    .ZN(_06260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14263_ (.A1(_04530_),
    .A2(_06015_),
    .ZN(_06261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14264_ (.A1(\filters.band[27] ),
    .A2(_04590_),
    .ZN(_06262_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14265_ (.A1(_06260_),
    .A2(_06261_),
    .A3(_06262_),
    .ZN(_06263_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14266_ (.A1(_04602_),
    .A2(_05802_),
    .A3(_06178_),
    .ZN(_06264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14267_ (.A1(_06176_),
    .A2(_06177_),
    .B(_06264_),
    .ZN(_06265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14268_ (.A1(_04728_),
    .A2(_05534_),
    .ZN(_06266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14269_ (.A1(_04251_),
    .A2(_05717_),
    .ZN(_06267_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14270_ (.A1(_06266_),
    .A2(_06267_),
    .Z(_06268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14271_ (.A1(_04261_),
    .A2(_05918_),
    .ZN(_06269_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14272_ (.A1(_06268_),
    .A2(_06269_),
    .ZN(_06270_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14273_ (.A1(_06265_),
    .A2(_06270_),
    .Z(_06271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14274_ (.A1(_06263_),
    .A2(_06271_),
    .Z(_06272_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14275_ (.A1(_06259_),
    .A2(_06272_),
    .Z(_06273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14276_ (.A1(_06256_),
    .A2(_06273_),
    .Z(_06274_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14277_ (.A1(_06253_),
    .A2(_06274_),
    .Z(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14278_ (.A1(_06217_),
    .A2(_06275_),
    .Z(_06276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14279_ (.I(_05586_),
    .Z(_06277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14280_ (.I(_06119_),
    .Z(_06278_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14281_ (.A1(_06277_),
    .A2(_06278_),
    .A3(_06121_),
    .ZN(_06279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14282_ (.A1(_06008_),
    .A2(_06112_),
    .A3(_06123_),
    .ZN(_06280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14283_ (.A1(_06279_),
    .A2(_06280_),
    .Z(_06281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14284_ (.A1(_06167_),
    .A2(_06182_),
    .ZN(_06282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14285_ (.A1(_06164_),
    .A2(_06183_),
    .B(_06282_),
    .ZN(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14286_ (.A1(_06169_),
    .A2(_06170_),
    .Z(_06284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14287_ (.I(_06034_),
    .Z(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14288_ (.A1(_04645_),
    .A2(_06285_),
    .A3(_06171_),
    .ZN(_06286_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14289_ (.A1(_06284_),
    .A2(_06286_),
    .Z(_06287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14290_ (.A1(_04674_),
    .A2(_06285_),
    .ZN(_06288_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14291_ (.A1(_06287_),
    .A2(_06288_),
    .ZN(_06289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14292_ (.A1(_04669_),
    .A2(_06278_),
    .ZN(_06290_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14293_ (.A1(_06289_),
    .A2(_06290_),
    .Z(_06291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14294_ (.A1(_06289_),
    .A2(_06290_),
    .ZN(_06292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14295_ (.A1(_06291_),
    .A2(_06292_),
    .ZN(_06293_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14296_ (.A1(_06283_),
    .A2(_06293_),
    .Z(_06294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14297_ (.A1(_06283_),
    .A2(_06293_),
    .ZN(_06295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14298_ (.A1(_06294_),
    .A2(_06295_),
    .ZN(_06296_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14299_ (.A1(_06281_),
    .A2(_06296_),
    .Z(_06297_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14300_ (.A1(_06276_),
    .A2(_06297_),
    .Z(_06298_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _14301_ (.A1(_06212_),
    .A2(_06215_),
    .A3(_06298_),
    .ZN(_06299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14302_ (.A1(_06111_),
    .A2(_06187_),
    .ZN(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _14303_ (.A1(_06108_),
    .A2(_06188_),
    .B(_06300_),
    .ZN(_06301_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14304_ (.A1(_06299_),
    .A2(_06301_),
    .Z(_06302_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14305_ (.I(_06193_),
    .ZN(_06303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14306_ (.A1(_06189_),
    .A2(_06192_),
    .ZN(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _14307_ (.I(_06304_),
    .ZN(_06305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14308_ (.A1(_06303_),
    .A2(_06200_),
    .B(_06305_),
    .ZN(_06306_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14309_ (.A1(_06306_),
    .A2(_06302_),
    .ZN(_06307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14310_ (.A1(_03347_),
    .A2(_05880_),
    .ZN(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _14311_ (.A1(_03349_),
    .A2(_06202_),
    .B(_06308_),
    .ZN(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14312_ (.A1(_06307_),
    .A2(_06309_),
    .Z(_06310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14313_ (.I(_06201_),
    .Z(_06311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14314_ (.A1(_06311_),
    .A2(_06204_),
    .ZN(_06312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14315_ (.A1(_06311_),
    .A2(_06204_),
    .ZN(_06313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14316_ (.A1(_06312_),
    .A2(_06208_),
    .B(_06313_),
    .ZN(_06314_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14317_ (.A1(_06310_),
    .A2(_06314_),
    .Z(_06315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14318_ (.A1(_06000_),
    .A2(_06315_),
    .ZN(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14319_ (.A1(_03349_),
    .A2(_06106_),
    .B(_06316_),
    .C(_06105_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14320_ (.I(_06307_),
    .Z(_06317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14321_ (.I(_06317_),
    .Z(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14322_ (.A1(_06318_),
    .A2(_06309_),
    .ZN(_06319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _14323_ (.A1(_06311_),
    .A2(_06204_),
    .B1(_06317_),
    .B2(_06309_),
    .ZN(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14324_ (.A1(_06205_),
    .A2(_06310_),
    .ZN(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _14325_ (.A1(_06319_),
    .A2(_06320_),
    .B1(_06321_),
    .B2(_06208_),
    .ZN(_06322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14326_ (.A1(_06193_),
    .A2(_06302_),
    .ZN(_06323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14327_ (.A1(_06194_),
    .A2(_06323_),
    .ZN(_06324_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14328_ (.A1(_06299_),
    .A2(_06301_),
    .Z(_06325_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _14329_ (.A1(_06305_),
    .A2(_06325_),
    .B1(_06323_),
    .B2(_06198_),
    .ZN(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14330_ (.A1(_06299_),
    .A2(_06301_),
    .ZN(_06327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _14331_ (.A1(_05904_),
    .A2(_06324_),
    .B(_06326_),
    .C(_06327_),
    .ZN(_06328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14332_ (.A1(_06281_),
    .A2(_06296_),
    .B(_06294_),
    .ZN(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14333_ (.A1(_06217_),
    .A2(_06275_),
    .ZN(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14334_ (.A1(_06276_),
    .A2(_06297_),
    .ZN(_06331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14335_ (.A1(_06330_),
    .A2(_06331_),
    .ZN(_06332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14336_ (.A1(_06220_),
    .A2(_06252_),
    .ZN(_06333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14337_ (.A1(_06253_),
    .A2(_06274_),
    .ZN(_06334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14338_ (.A1(_06333_),
    .A2(_06334_),
    .ZN(_06335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14339_ (.A1(_06224_),
    .A2(_06238_),
    .ZN(_06336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14340_ (.A1(_06239_),
    .A2(_06251_),
    .ZN(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14341_ (.A1(_06336_),
    .A2(_06337_),
    .ZN(_06338_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14342_ (.A1(_06233_),
    .A2(_06237_),
    .Z(_06339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14343_ (.A1(_06227_),
    .A2(_06232_),
    .B(_06339_),
    .ZN(_06340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14344_ (.A1(_06228_),
    .A2(_06229_),
    .ZN(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14345_ (.A1(_06230_),
    .A2(_06231_),
    .ZN(_06342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14346_ (.A1(_06341_),
    .A2(_06342_),
    .ZN(_06343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14347_ (.A1(_05496_),
    .A2(_05651_),
    .ZN(_06344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14348_ (.A1(_04889_),
    .A2(_05516_),
    .ZN(_06345_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14349_ (.A1(_06344_),
    .A2(_06345_),
    .ZN(_06346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14350_ (.A1(_04850_),
    .A2(_05076_),
    .ZN(_06347_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14351_ (.A1(_06346_),
    .A2(_06347_),
    .ZN(_06348_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14352_ (.A1(_06343_),
    .A2(_06348_),
    .ZN(_06349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14353_ (.A1(_05959_),
    .A2(_05119_),
    .ZN(_06350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14354_ (.A1(_05857_),
    .A2(_05306_),
    .ZN(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14355_ (.A1(_04475_),
    .A2(_05396_),
    .ZN(_06352_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14356_ (.A1(_06350_),
    .A2(_06351_),
    .A3(_06352_),
    .Z(_06353_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14357_ (.A1(_06349_),
    .A2(_06353_),
    .Z(_06354_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14358_ (.A1(_06340_),
    .A2(_06354_),
    .Z(_06355_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14359_ (.A1(_04386_),
    .A2(_05596_),
    .A3(_06248_),
    .ZN(_06356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14360_ (.A1(_06246_),
    .A2(_06247_),
    .B(_06356_),
    .ZN(_06357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14361_ (.A1(_06234_),
    .A2(_06235_),
    .ZN(_06358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14362_ (.A1(_06234_),
    .A2(_06235_),
    .ZN(_06359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14363_ (.A1(_06358_),
    .A2(_06236_),
    .B(_06359_),
    .ZN(_06360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14364_ (.A1(_04355_),
    .A2(_05699_),
    .ZN(_06361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14365_ (.A1(_04407_),
    .A2(_05947_),
    .ZN(_06362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14366_ (.A1(_04477_),
    .A2(_05529_),
    .ZN(_06363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14367_ (.A1(_06362_),
    .A2(_06363_),
    .Z(_06364_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14368_ (.A1(_06361_),
    .A2(_06364_),
    .ZN(_06365_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14369_ (.A1(_06360_),
    .A2(_06365_),
    .Z(_06366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14370_ (.I(_06366_),
    .ZN(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14371_ (.A1(_06357_),
    .A2(_06367_),
    .Z(_06368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14372_ (.A1(_06355_),
    .A2(_06368_),
    .Z(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14373_ (.A1(_06338_),
    .A2(_06369_),
    .Z(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14374_ (.A1(_06265_),
    .A2(_06270_),
    .ZN(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14375_ (.A1(_06263_),
    .A2(_06271_),
    .ZN(_06372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14376_ (.A1(_06371_),
    .A2(_06372_),
    .ZN(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14377_ (.A1(_06244_),
    .A2(_06249_),
    .ZN(_06374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14378_ (.A1(_06242_),
    .A2(_06250_),
    .ZN(_06375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14379_ (.A1(_06374_),
    .A2(_06375_),
    .ZN(_06376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14380_ (.A1(\filters.band[27] ),
    .A2(_04606_),
    .ZN(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14381_ (.A1(_04628_),
    .A2(_06119_),
    .ZN(_06378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14382_ (.I(\filters.band[28] ),
    .Z(_06379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14383_ (.A1(_06379_),
    .A2(_04627_),
    .ZN(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14384_ (.A1(_06377_),
    .A2(_06378_),
    .A3(_06380_),
    .ZN(_06381_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14385_ (.A1(_04603_),
    .A2(_05921_),
    .A3(_06268_),
    .ZN(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14386_ (.A1(_06266_),
    .A2(_06267_),
    .B(_06382_),
    .ZN(_06383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14387_ (.A1(_04602_),
    .A2(_06015_),
    .ZN(_06384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14388_ (.I(_04271_),
    .Z(_06385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14389_ (.A1(_06385_),
    .A2(_05717_),
    .ZN(_06386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14390_ (.A1(_05540_),
    .A2(_05821_),
    .ZN(_06387_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14391_ (.A1(_06386_),
    .A2(_06387_),
    .Z(_06388_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14392_ (.A1(_06384_),
    .A2(_06388_),
    .ZN(_06389_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14393_ (.A1(_06383_),
    .A2(_06389_),
    .Z(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14394_ (.A1(_06381_),
    .A2(_06390_),
    .Z(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14395_ (.A1(_06376_),
    .A2(_06391_),
    .Z(_06392_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14396_ (.A1(_06373_),
    .A2(_06392_),
    .Z(_06393_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14397_ (.A1(_06370_),
    .A2(_06393_),
    .Z(_06394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14398_ (.A1(_06335_),
    .A2(_06394_),
    .Z(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14399_ (.A1(_06287_),
    .A2(_06288_),
    .B(_06291_),
    .ZN(_06396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14400_ (.A1(_06259_),
    .A2(_06272_),
    .ZN(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14401_ (.A1(_06256_),
    .A2(_06273_),
    .ZN(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14402_ (.A1(_06397_),
    .A2(_06398_),
    .ZN(_06399_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14403_ (.A1(_06261_),
    .A2(_06262_),
    .Z(_06400_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14404_ (.A1(_06261_),
    .A2(_06262_),
    .Z(_06401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14405_ (.A1(_06260_),
    .A2(_06400_),
    .B(_06401_),
    .ZN(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14406_ (.I(\filters.band[26] ),
    .Z(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14407_ (.A1(_06403_),
    .A2(_04661_),
    .ZN(_06404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14408_ (.A1(_06402_),
    .A2(_06404_),
    .ZN(_06405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14409_ (.I(_06285_),
    .Z(_06406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14410_ (.A1(_05589_),
    .A2(_06406_),
    .ZN(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14411_ (.A1(_06405_),
    .A2(_06407_),
    .ZN(_06408_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14412_ (.A1(_06399_),
    .A2(_06408_),
    .Z(_06409_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14413_ (.A1(_06396_),
    .A2(_06409_),
    .Z(_06410_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14414_ (.A1(_06395_),
    .A2(_06410_),
    .Z(_06411_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14415_ (.A1(_06332_),
    .A2(_06411_),
    .Z(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14416_ (.A1(_06329_),
    .A2(_06412_),
    .Z(_06413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14417_ (.A1(_06215_),
    .A2(_06298_),
    .ZN(_06414_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14418_ (.A1(_06215_),
    .A2(_06298_),
    .Z(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14419_ (.A1(_06212_),
    .A2(_06414_),
    .A3(_06415_),
    .ZN(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _14420_ (.A1(_06414_),
    .A2(_06416_),
    .ZN(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14421_ (.A1(_06413_),
    .A2(_06417_),
    .ZN(_06418_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14422_ (.A1(_06328_),
    .A2(_06418_),
    .ZN(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14423_ (.I(_05880_),
    .Z(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14424_ (.A1(_03362_),
    .A2(_03223_),
    .ZN(_06421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14425_ (.A1(_03363_),
    .A2(_06420_),
    .B(_06421_),
    .ZN(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14426_ (.A1(_06419_),
    .A2(_06422_),
    .Z(_06423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14427_ (.A1(_06322_),
    .A2(_06423_),
    .Z(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14428_ (.A1(_06000_),
    .A2(_06424_),
    .ZN(_06425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14429_ (.A1(_03363_),
    .A2(_06106_),
    .B(_06425_),
    .C(_06105_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14430_ (.I(_05569_),
    .Z(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14431_ (.A1(_06399_),
    .A2(_06408_),
    .ZN(_06427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14432_ (.A1(_06396_),
    .A2(_06409_),
    .ZN(_06428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14433_ (.A1(_06427_),
    .A2(_06428_),
    .ZN(_06429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14434_ (.A1(_06335_),
    .A2(_06394_),
    .ZN(_06430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14435_ (.A1(_06395_),
    .A2(_06410_),
    .ZN(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14436_ (.A1(_06430_),
    .A2(_06431_),
    .ZN(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14437_ (.A1(_06338_),
    .A2(_06369_),
    .ZN(_06433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14438_ (.A1(_06370_),
    .A2(_06393_),
    .ZN(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14439_ (.A1(_06433_),
    .A2(_06434_),
    .ZN(_06435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14440_ (.A1(_06340_),
    .A2(_06354_),
    .ZN(_06436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14441_ (.A1(_06355_),
    .A2(_06368_),
    .ZN(_06437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14442_ (.A1(_06436_),
    .A2(_06437_),
    .ZN(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14443_ (.A1(_06343_),
    .A2(_06348_),
    .Z(_06439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14444_ (.A1(_06349_),
    .A2(_06353_),
    .B(_06439_),
    .ZN(_06440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14445_ (.A1(_06344_),
    .A2(_06345_),
    .ZN(_06441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14446_ (.A1(_06346_),
    .A2(_06347_),
    .ZN(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14447_ (.A1(_06441_),
    .A2(_06442_),
    .ZN(_06443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14448_ (.A1(_05617_),
    .A2(_05652_),
    .ZN(_06444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14449_ (.A1(_04952_),
    .A2(_05650_),
    .ZN(_06445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14450_ (.A1(_04851_),
    .A2(_05119_),
    .ZN(_06446_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14451_ (.A1(_06444_),
    .A2(_06445_),
    .A3(_06446_),
    .Z(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14452_ (.A1(_06443_),
    .A2(_06447_),
    .Z(_06448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14453_ (.A1(_05751_),
    .A2(_05305_),
    .ZN(_06449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14454_ (.A1(_04837_),
    .A2(_05395_),
    .ZN(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14455_ (.A1(_06449_),
    .A2(_06450_),
    .Z(_06451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14456_ (.A1(_04475_),
    .A2(_05474_),
    .ZN(_06452_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14457_ (.A1(_06451_),
    .A2(_06452_),
    .ZN(_06453_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14458_ (.A1(_06448_),
    .A2(_06453_),
    .Z(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14459_ (.A1(_06440_),
    .A2(_06454_),
    .Z(_06455_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14460_ (.A1(_06362_),
    .A2(_06363_),
    .Z(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14461_ (.I(_04386_),
    .Z(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14462_ (.A1(_06457_),
    .A2(_05700_),
    .A3(_06364_),
    .ZN(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14463_ (.A1(_06456_),
    .A2(_06458_),
    .Z(_06459_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14464_ (.A1(_06350_),
    .A2(_06351_),
    .Z(_06460_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14465_ (.A1(_06350_),
    .A2(_06351_),
    .Z(_06461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14466_ (.A1(_06460_),
    .A2(_06352_),
    .B(_06461_),
    .ZN(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14467_ (.A1(_04386_),
    .A2(_05802_),
    .ZN(_06463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14468_ (.A1(_04481_),
    .A2(_05529_),
    .ZN(_06464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14469_ (.A1(_04347_),
    .A2(_05699_),
    .ZN(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14470_ (.A1(_06464_),
    .A2(_06465_),
    .Z(_06466_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14471_ (.A1(_06463_),
    .A2(_06466_),
    .ZN(_06467_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14472_ (.A1(_06462_),
    .A2(_06467_),
    .ZN(_06468_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14473_ (.A1(_06459_),
    .A2(_06468_),
    .Z(_06469_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14474_ (.A1(_06455_),
    .A2(_06469_),
    .Z(_06470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14475_ (.A1(_06438_),
    .A2(_06470_),
    .Z(_06471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14476_ (.A1(_06383_),
    .A2(_06389_),
    .ZN(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14477_ (.A1(_06381_),
    .A2(_06390_),
    .ZN(_06473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14478_ (.A1(_06472_),
    .A2(_06473_),
    .ZN(_06474_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14479_ (.I(_06365_),
    .ZN(_06475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14480_ (.A1(_06357_),
    .A2(_06367_),
    .ZN(_06476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14481_ (.A1(_06360_),
    .A2(_06475_),
    .B(_06476_),
    .ZN(_06477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14482_ (.A1(\filters.band[28] ),
    .A2(_04625_),
    .ZN(_06478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14483_ (.A1(_04628_),
    .A2(_06034_),
    .ZN(_06479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14484_ (.A1(\filters.band[29] ),
    .A2(_04646_),
    .ZN(_06480_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14485_ (.A1(_06478_),
    .A2(_06479_),
    .A3(_06480_),
    .ZN(_06481_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14486_ (.A1(_04603_),
    .A2(_06016_),
    .A3(_06388_),
    .ZN(_06482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14487_ (.A1(_06386_),
    .A2(_06387_),
    .B(_06482_),
    .ZN(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14488_ (.A1(_04602_),
    .A2(_06031_),
    .ZN(_06484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14489_ (.A1(_06385_),
    .A2(_05821_),
    .ZN(_06485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14490_ (.A1(_04252_),
    .A2(_05824_),
    .ZN(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14491_ (.A1(_06485_),
    .A2(_06486_),
    .Z(_06487_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14492_ (.A1(_06484_),
    .A2(_06487_),
    .ZN(_06488_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14493_ (.A1(_06483_),
    .A2(_06488_),
    .Z(_06489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14494_ (.A1(_06481_),
    .A2(_06489_),
    .Z(_06490_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14495_ (.A1(_06477_),
    .A2(_06490_),
    .Z(_06491_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14496_ (.A1(_06474_),
    .A2(_06491_),
    .Z(_06492_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14497_ (.A1(_06471_),
    .A2(_06492_),
    .Z(_06493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14498_ (.A1(_06435_),
    .A2(_06493_),
    .Z(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14499_ (.I(_06403_),
    .Z(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14500_ (.I(_06277_),
    .Z(_06496_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14501_ (.A1(_06495_),
    .A2(_06496_),
    .A3(_06402_),
    .ZN(_06497_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14502_ (.A1(_06008_),
    .A2(_06406_),
    .A3(_06405_),
    .ZN(_06498_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14503_ (.A1(_06497_),
    .A2(_06498_),
    .Z(_06499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14504_ (.A1(_06376_),
    .A2(_06391_),
    .ZN(_06500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14505_ (.A1(_06373_),
    .A2(_06392_),
    .ZN(_06501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14506_ (.A1(_06500_),
    .A2(_06501_),
    .ZN(_06502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14507_ (.A1(_06403_),
    .A2(_05589_),
    .ZN(_06503_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14508_ (.A1(_06378_),
    .A2(_06380_),
    .Z(_06504_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14509_ (.A1(_06378_),
    .A2(_06380_),
    .Z(_06505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14510_ (.A1(_06377_),
    .A2(_06504_),
    .B(_06505_),
    .ZN(_06506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14511_ (.I(\filters.band[27] ),
    .Z(_06507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14512_ (.A1(_06507_),
    .A2(_05586_),
    .ZN(_06508_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14513_ (.A1(_06503_),
    .A2(_06506_),
    .A3(_06508_),
    .Z(_06509_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14514_ (.A1(_06502_),
    .A2(_06509_),
    .ZN(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14515_ (.A1(_06499_),
    .A2(_06510_),
    .Z(_06511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14516_ (.A1(_06494_),
    .A2(_06511_),
    .Z(_06512_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14517_ (.A1(_06429_),
    .A2(_06432_),
    .A3(_06512_),
    .ZN(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14518_ (.A1(_06332_),
    .A2(_06411_),
    .ZN(_06514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14519_ (.A1(_06329_),
    .A2(_06412_),
    .ZN(_06515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14520_ (.A1(_06514_),
    .A2(_06515_),
    .ZN(_06516_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14521_ (.A1(_06513_),
    .A2(_06516_),
    .Z(_06517_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14522_ (.A1(_06413_),
    .A2(_06417_),
    .Z(_06518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14523_ (.I(_06518_),
    .ZN(_06519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14524_ (.A1(_06328_),
    .A2(_06418_),
    .B(_06519_),
    .ZN(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14525_ (.A1(_06517_),
    .A2(_06520_),
    .Z(_06521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14526_ (.I(_06521_),
    .Z(_06522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14527_ (.A1(_03376_),
    .A2(_06202_),
    .ZN(_06523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14528_ (.A1(_03382_),
    .A2(_03380_),
    .B(_06523_),
    .ZN(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14529_ (.A1(_06522_),
    .A2(_06524_),
    .Z(_06525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14530_ (.A1(_06419_),
    .A2(_06422_),
    .ZN(_06526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14531_ (.A1(_06322_),
    .A2(_06423_),
    .ZN(_06527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14532_ (.A1(_06526_),
    .A2(_06527_),
    .ZN(_06528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14533_ (.A1(_06525_),
    .A2(_06528_),
    .Z(_06529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14534_ (.A1(_06426_),
    .A2(_06529_),
    .ZN(_06530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14535_ (.I(_01827_),
    .Z(_06531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14536_ (.A1(_03382_),
    .A2(_06106_),
    .B(_06530_),
    .C(_06531_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14537_ (.I(_05570_),
    .Z(_06532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14538_ (.A1(_06514_),
    .A2(_06515_),
    .B(_06513_),
    .ZN(_06533_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14539_ (.A1(_06514_),
    .A2(_06515_),
    .A3(_06513_),
    .ZN(_06534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14540_ (.A1(_06518_),
    .A2(_06533_),
    .B(_06534_),
    .ZN(_06535_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _14541_ (.A1(_06328_),
    .A2(_06418_),
    .A3(_06517_),
    .B(_06535_),
    .ZN(_06536_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14542_ (.A1(_06432_),
    .A2(_06512_),
    .Z(_06537_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14543_ (.A1(_06432_),
    .A2(_06512_),
    .Z(_06538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14544_ (.A1(_06429_),
    .A2(_06537_),
    .B(_06538_),
    .ZN(_06539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14545_ (.A1(_06502_),
    .A2(_06509_),
    .ZN(_06540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14546_ (.A1(_06499_),
    .A2(_06510_),
    .B(_06540_),
    .ZN(_06541_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14547_ (.A1(_06435_),
    .A2(_06493_),
    .Z(_06542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14548_ (.A1(_06494_),
    .A2(_06511_),
    .B(_06542_),
    .ZN(_06543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14549_ (.I(_06507_),
    .Z(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14550_ (.A1(_06544_),
    .A2(_06277_),
    .B(_06506_),
    .ZN(_06545_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14551_ (.A1(_06507_),
    .A2(_06277_),
    .A3(_06506_),
    .ZN(_06546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14552_ (.A1(_06503_),
    .A2(_06545_),
    .B(_06546_),
    .ZN(_06547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14553_ (.A1(_06477_),
    .A2(_06490_),
    .ZN(_06548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14554_ (.A1(_06474_),
    .A2(_06491_),
    .ZN(_06549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14555_ (.A1(_06548_),
    .A2(_06549_),
    .ZN(_06550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14556_ (.A1(_06507_),
    .A2(_04660_),
    .ZN(_06551_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14557_ (.A1(_06479_),
    .A2(_06480_),
    .Z(_06552_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14558_ (.A1(_06479_),
    .A2(_06480_),
    .Z(_06553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14559_ (.A1(_06478_),
    .A2(_06552_),
    .B(_06553_),
    .ZN(_06554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14560_ (.A1(_06379_),
    .A2(_04697_),
    .ZN(_06555_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14561_ (.A1(_06551_),
    .A2(_06554_),
    .A3(_06555_),
    .Z(_06556_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14562_ (.A1(_06550_),
    .A2(_06556_),
    .Z(_06557_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14563_ (.A1(_06547_),
    .A2(_06557_),
    .ZN(_06558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14564_ (.A1(_06438_),
    .A2(_06470_),
    .ZN(_06559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14565_ (.A1(_06471_),
    .A2(_06492_),
    .ZN(_06560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14566_ (.A1(_06559_),
    .A2(_06560_),
    .ZN(_06561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14567_ (.A1(_06483_),
    .A2(_06488_),
    .ZN(_06562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14568_ (.A1(_06481_),
    .A2(_06489_),
    .ZN(_06563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14569_ (.A1(_06562_),
    .A2(_06563_),
    .ZN(_06564_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14570_ (.I(_06564_),
    .ZN(_06565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14571_ (.A1(_06462_),
    .A2(_06467_),
    .ZN(_06566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14572_ (.A1(_06459_),
    .A2(_06468_),
    .B(_06566_),
    .ZN(_06567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14573_ (.I(\filters.band[29] ),
    .Z(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14574_ (.A1(_06568_),
    .A2(_04645_),
    .ZN(_06569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14575_ (.A1(_06403_),
    .A2(_04629_),
    .ZN(_06570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14576_ (.A1(\filters.band[30] ),
    .A2(_04627_),
    .ZN(_06571_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14577_ (.A1(_06570_),
    .A2(_06571_),
    .Z(_06572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14578_ (.A1(_06570_),
    .A2(_06571_),
    .ZN(_06573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14579_ (.A1(_06572_),
    .A2(_06573_),
    .ZN(_06574_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14580_ (.A1(_06569_),
    .A2(_06574_),
    .Z(_06575_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14581_ (.A1(_04604_),
    .A2(_06278_),
    .A3(_06487_),
    .ZN(_06576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14582_ (.A1(_06485_),
    .A2(_06486_),
    .B(_06576_),
    .ZN(_06577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14583_ (.A1(_04603_),
    .A2(_06285_),
    .ZN(_06578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14584_ (.A1(_06385_),
    .A2(_06015_),
    .ZN(_06579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14585_ (.A1(_04252_),
    .A2(_06031_),
    .ZN(_06580_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14586_ (.A1(_06579_),
    .A2(_06580_),
    .Z(_06581_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14587_ (.A1(_06578_),
    .A2(_06581_),
    .ZN(_06582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14588_ (.A1(_06577_),
    .A2(_06582_),
    .Z(_06583_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14589_ (.A1(_06575_),
    .A2(_06583_),
    .Z(_06584_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14590_ (.A1(_06565_),
    .A2(_06567_),
    .A3(_06584_),
    .Z(_06585_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14591_ (.A1(_06440_),
    .A2(_06454_),
    .Z(_06586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14592_ (.A1(_06455_),
    .A2(_06469_),
    .B(_06586_),
    .ZN(_06587_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14593_ (.A1(_06464_),
    .A2(_06465_),
    .Z(_06588_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14594_ (.A1(_06457_),
    .A2(_05803_),
    .A3(_06466_),
    .ZN(_06589_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14595_ (.A1(_06588_),
    .A2(_06589_),
    .Z(_06590_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14596_ (.A1(_05713_),
    .A2(_05475_),
    .A3(_06451_),
    .ZN(_06591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14597_ (.A1(_06449_),
    .A2(_06450_),
    .B(_06591_),
    .ZN(_06592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14598_ (.A1(_04355_),
    .A2(_05918_),
    .ZN(_06593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14599_ (.A1(_04481_),
    .A2(_05699_),
    .ZN(_06594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14600_ (.A1(_04347_),
    .A2(_05802_),
    .ZN(_06595_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14601_ (.A1(_06594_),
    .A2(_06595_),
    .Z(_06596_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14602_ (.A1(_06593_),
    .A2(_06596_),
    .ZN(_06597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14603_ (.A1(_06592_),
    .A2(_06597_),
    .Z(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14604_ (.A1(_06590_),
    .A2(_06598_),
    .Z(_06599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14605_ (.A1(_06443_),
    .A2(_06447_),
    .ZN(_06600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14606_ (.A1(_06448_),
    .A2(_06453_),
    .B(_06600_),
    .ZN(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14607_ (.A1(_04474_),
    .A2(_05530_),
    .ZN(_06602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14608_ (.A1(_05959_),
    .A2(_05396_),
    .ZN(_06603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14609_ (.A1(_05857_),
    .A2(_05474_),
    .ZN(_06604_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14610_ (.A1(_06602_),
    .A2(_06603_),
    .A3(_06604_),
    .ZN(_06605_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14611_ (.A1(_06444_),
    .A2(_06445_),
    .Z(_06606_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14612_ (.A1(_06444_),
    .A2(_06445_),
    .Z(_06607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14613_ (.A1(_06606_),
    .A2(_06446_),
    .B(_06607_),
    .ZN(_06608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14614_ (.A1(_04851_),
    .A2(_05306_),
    .ZN(_06609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14615_ (.A1(_05077_),
    .A2(_05652_),
    .ZN(_06610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14616_ (.A1(_05650_),
    .A2(_05120_),
    .ZN(_06611_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14617_ (.A1(_06609_),
    .A2(_06610_),
    .A3(_06611_),
    .ZN(_06612_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14618_ (.A1(_06608_),
    .A2(_06612_),
    .Z(_06613_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14619_ (.A1(_06601_),
    .A2(_06605_),
    .A3(_06613_),
    .Z(_06614_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14620_ (.A1(_06599_),
    .A2(_06614_),
    .ZN(_06615_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14621_ (.A1(_06587_),
    .A2(_06615_),
    .Z(_06616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14622_ (.A1(_06587_),
    .A2(_06615_),
    .ZN(_06617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14623_ (.A1(_06616_),
    .A2(_06617_),
    .ZN(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14624_ (.A1(_06618_),
    .A2(_06585_),
    .Z(_06619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14625_ (.A1(_06561_),
    .A2(_06619_),
    .Z(_06620_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14626_ (.A1(_06558_),
    .A2(_06620_),
    .ZN(_06621_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14627_ (.A1(_06543_),
    .A2(_06621_),
    .ZN(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14628_ (.A1(_06541_),
    .A2(_06622_),
    .ZN(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14629_ (.A1(_06539_),
    .A2(_06623_),
    .Z(_06624_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14630_ (.A1(net30),
    .A2(_06624_),
    .ZN(_06625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14631_ (.A1(\filters.low[10] ),
    .A2(_03379_),
    .ZN(_06626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14632_ (.A1(_03398_),
    .A2(_06092_),
    .B(_06626_),
    .ZN(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14633_ (.A1(_06625_),
    .A2(_06627_),
    .ZN(_06628_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14634_ (.A1(_06423_),
    .A2(_06525_),
    .Z(_06629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14635_ (.A1(_06522_),
    .A2(_06524_),
    .ZN(_06630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14636_ (.A1(_06522_),
    .A2(_06524_),
    .ZN(_06631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14637_ (.A1(_06526_),
    .A2(_06630_),
    .B(_06631_),
    .ZN(_06632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14638_ (.A1(_06322_),
    .A2(_06629_),
    .B(_06632_),
    .ZN(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14639_ (.A1(net32),
    .A2(_06633_),
    .Z(_06634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14640_ (.A1(_06426_),
    .A2(_06634_),
    .ZN(_06635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14641_ (.A1(_03398_),
    .A2(_06532_),
    .B(_06635_),
    .C(_06531_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14642_ (.I(_06543_),
    .ZN(_06636_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14643_ (.A1(_06636_),
    .A2(_06621_),
    .Z(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14644_ (.A1(_06541_),
    .A2(_06622_),
    .B(_06637_),
    .ZN(_06638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14645_ (.I(_06379_),
    .Z(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14646_ (.A1(_06639_),
    .A2(_06496_),
    .B(_06554_),
    .ZN(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14647_ (.A1(_06639_),
    .A2(_06496_),
    .A3(_06554_),
    .ZN(_06641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14648_ (.A1(_06551_),
    .A2(_06640_),
    .B(_06641_),
    .ZN(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14649_ (.A1(_06385_),
    .A2(_06278_),
    .ZN(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14650_ (.A1(_06577_),
    .A2(_06582_),
    .ZN(_06644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14651_ (.A1(_06575_),
    .A2(_06583_),
    .ZN(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14652_ (.A1(_06644_),
    .A2(_06645_),
    .ZN(_06646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14653_ (.A1(\filters.band[31] ),
    .A2(_04665_),
    .ZN(_06647_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14654_ (.A1(_06643_),
    .A2(_06646_),
    .A3(_06647_),
    .Z(_06648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14655_ (.A1(_06495_),
    .A2(_04604_),
    .ZN(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14656_ (.A1(_04604_),
    .A2(_06406_),
    .A3(_06581_),
    .ZN(_06650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14657_ (.A1(_06579_),
    .A2(_06580_),
    .B(_06650_),
    .ZN(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14658_ (.A1(_06585_),
    .A2(_06618_),
    .B(_06616_),
    .ZN(_06652_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14659_ (.A1(_06649_),
    .A2(_06651_),
    .A3(_06652_),
    .Z(_06653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14660_ (.A1(_06544_),
    .A2(_04629_),
    .ZN(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14661_ (.I(_06598_),
    .ZN(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14662_ (.A1(_06592_),
    .A2(_06597_),
    .ZN(_06656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14663_ (.A1(_06590_),
    .A2(_06655_),
    .B(_06656_),
    .ZN(_06657_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14664_ (.A1(_06610_),
    .A2(_06611_),
    .Z(_06658_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14665_ (.A1(_06610_),
    .A2(_06611_),
    .Z(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14666_ (.A1(_06609_),
    .A2(_06658_),
    .B(_06659_),
    .ZN(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14667_ (.A1(_05713_),
    .A2(_05794_),
    .ZN(_06661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14668_ (.A1(_05650_),
    .A2(_05307_),
    .ZN(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14669_ (.A1(_05959_),
    .A2(_05587_),
    .ZN(_06663_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14670_ (.A1(_06603_),
    .A2(_06604_),
    .Z(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14671_ (.A1(_06603_),
    .A2(_06604_),
    .Z(_06665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14672_ (.A1(_06602_),
    .A2(_06664_),
    .B(_06665_),
    .ZN(_06666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14673_ (.A1(_04347_),
    .A2(_06006_),
    .ZN(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14674_ (.A1(_06663_),
    .A2(_06666_),
    .A3(_06667_),
    .Z(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14675_ (.A1(_06661_),
    .A2(_06662_),
    .A3(_06668_),
    .Z(_06669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14676_ (.A1(_04252_),
    .A2(_06406_),
    .ZN(_06670_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14677_ (.A1(_06660_),
    .A2(_06669_),
    .A3(_06670_),
    .Z(_06671_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14678_ (.A1(_06654_),
    .A2(_06657_),
    .A3(_06671_),
    .Z(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14679_ (.A1(_06648_),
    .A2(_06653_),
    .A3(_06672_),
    .Z(_06673_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14680_ (.A1(_06638_),
    .A2(_06642_),
    .A3(_06673_),
    .Z(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14681_ (.A1(_06569_),
    .A2(_06574_),
    .B(_06572_),
    .ZN(_06675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14682_ (.A1(_04481_),
    .A2(_05910_),
    .ZN(_06676_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14683_ (.A1(_06457_),
    .A2(_06006_),
    .A3(_06596_),
    .ZN(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14684_ (.A1(_06594_),
    .A2(_06595_),
    .B(_06677_),
    .ZN(_06678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14685_ (.A1(\filters.band[30] ),
    .A2(_04662_),
    .ZN(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14686_ (.A1(_06676_),
    .A2(_06678_),
    .A3(_06679_),
    .Z(_06680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14687_ (.A1(_06457_),
    .A2(_06112_),
    .ZN(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14688_ (.A1(_06605_),
    .A2(_06613_),
    .Z(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14689_ (.A1(_06605_),
    .A2(_06613_),
    .ZN(_06683_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _14690_ (.A1(_06601_),
    .A2(_06682_),
    .A3(_06683_),
    .B1(_06614_),
    .B2(_06599_),
    .ZN(_06684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14691_ (.A1(_06608_),
    .A2(_06612_),
    .ZN(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14692_ (.A1(_06605_),
    .A2(_06613_),
    .ZN(_06686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14693_ (.A1(_06685_),
    .A2(_06686_),
    .ZN(_06687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14694_ (.A1(_04851_),
    .A2(_05399_),
    .ZN(_06688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14695_ (.A1(_05294_),
    .A2(_05652_),
    .ZN(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14696_ (.A1(_05857_),
    .A2(_05691_),
    .ZN(_06690_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14697_ (.A1(_06688_),
    .A2(_06689_),
    .A3(_06690_),
    .Z(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14698_ (.A1(_06687_),
    .A2(_06691_),
    .Z(_06692_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14699_ (.A1(_06681_),
    .A2(_06684_),
    .A3(_06692_),
    .Z(_06693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14700_ (.A1(_06568_),
    .A2(_06496_),
    .ZN(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14701_ (.A1(_06680_),
    .A2(_06693_),
    .A3(_06694_),
    .Z(_06695_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14702_ (.I(_06620_),
    .ZN(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14703_ (.A1(_06561_),
    .A2(_06619_),
    .ZN(_06697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14704_ (.A1(_06558_),
    .A2(_06696_),
    .B(_06697_),
    .ZN(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14705_ (.A1(_06567_),
    .A2(_06584_),
    .ZN(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14706_ (.A1(_06567_),
    .A2(_06584_),
    .ZN(_06700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14707_ (.A1(_06565_),
    .A2(_06699_),
    .B(_06700_),
    .ZN(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14708_ (.A1(_06550_),
    .A2(_06556_),
    .ZN(_06702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14709_ (.A1(_06547_),
    .A2(_06557_),
    .ZN(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14710_ (.A1(_06702_),
    .A2(_06703_),
    .ZN(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14711_ (.A1(_06701_),
    .A2(_06704_),
    .Z(_06705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14712_ (.A1(_06379_),
    .A2(_06008_),
    .ZN(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14713_ (.A1(_06698_),
    .A2(_06705_),
    .A3(_06706_),
    .Z(_06707_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _14714_ (.A1(_06675_),
    .A2(_06695_),
    .A3(_06707_),
    .Z(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14715_ (.A1(_06539_),
    .A2(_06623_),
    .ZN(_06709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14716_ (.A1(_06536_),
    .A2(_06624_),
    .B(_06709_),
    .ZN(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _14717_ (.A1(_06674_),
    .A2(_06708_),
    .A3(_06710_),
    .Z(_06711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14718_ (.I(_06711_),
    .Z(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14719_ (.A1(_03413_),
    .A2(_03223_),
    .ZN(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14720_ (.A1(_03414_),
    .A2(_03380_),
    .B(_06713_),
    .ZN(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14721_ (.A1(_06712_),
    .A2(_06714_),
    .ZN(_06715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14722_ (.A1(_06625_),
    .A2(_06627_),
    .ZN(_06716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14723_ (.A1(net32),
    .A2(_06633_),
    .B(_06716_),
    .ZN(_06717_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14724_ (.A1(_06715_),
    .A2(_06717_),
    .Z(_06718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14725_ (.A1(\filters.band[11] ),
    .A2(_05567_),
    .B(_03753_),
    .ZN(_06719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14726_ (.A1(_04189_),
    .A2(_06718_),
    .B(_06719_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14727_ (.A1(_06423_),
    .A2(_06525_),
    .ZN(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _14728_ (.A1(_06628_),
    .A2(_06720_),
    .A3(_06715_),
    .ZN(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14729_ (.I(_06628_),
    .ZN(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _14730_ (.I(_06711_),
    .Z(_06723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _14731_ (.I(_06723_),
    .Z(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14732_ (.A1(_06724_),
    .A2(_06714_),
    .ZN(_06725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _14733_ (.I(_06723_),
    .Z(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _14734_ (.A1(_06726_),
    .A2(_06714_),
    .Z(_06727_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _14735_ (.A1(_06722_),
    .A2(_06632_),
    .A3(_06725_),
    .A4(_06727_),
    .Z(_06728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14736_ (.I(_06723_),
    .Z(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14737_ (.A1(_06729_),
    .A2(_06714_),
    .ZN(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14738_ (.A1(_06716_),
    .A2(_06730_),
    .B(_06725_),
    .ZN(_06731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _14739_ (.A1(_06322_),
    .A2(_06721_),
    .B(_06728_),
    .C(_06731_),
    .ZN(_06732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14740_ (.I(_06092_),
    .Z(_06733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14741_ (.A1(_03424_),
    .A2(_06420_),
    .ZN(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _14742_ (.A1(_03425_),
    .A2(_06733_),
    .B(_06734_),
    .ZN(_06735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14743_ (.A1(_06712_),
    .A2(_06735_),
    .Z(_06736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14744_ (.A1(_06732_),
    .A2(_06736_),
    .Z(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14745_ (.I(_03674_),
    .Z(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14746_ (.I(_06738_),
    .Z(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14747_ (.A1(\filters.band[12] ),
    .A2(_05567_),
    .B(_06739_),
    .ZN(_06740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14748_ (.A1(_04189_),
    .A2(_06737_),
    .B(_06740_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14749_ (.I(_06726_),
    .Z(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14750_ (.I(_06741_),
    .Z(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14751_ (.I(_06742_),
    .Z(_06743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14752_ (.I(_06743_),
    .Z(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14753_ (.I(_06744_),
    .Z(_06745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14754_ (.A1(_06745_),
    .A2(_06735_),
    .ZN(_06746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14755_ (.I(_06744_),
    .Z(_06747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14756_ (.A1(_06747_),
    .A2(_06735_),
    .ZN(_06748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14757_ (.A1(_06732_),
    .A2(_06746_),
    .B(_06748_),
    .ZN(_06749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14758_ (.A1(_03441_),
    .A2(_06733_),
    .ZN(_06750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14759_ (.A1(_03442_),
    .A2(_03224_),
    .B(_06750_),
    .ZN(_06751_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14760_ (.A1(_06712_),
    .A2(_06751_),
    .Z(_06752_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14761_ (.A1(_06749_),
    .A2(_06752_),
    .Z(_06753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14762_ (.A1(_06426_),
    .A2(_06753_),
    .ZN(_06754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14763_ (.A1(_03442_),
    .A2(_06532_),
    .B(_06754_),
    .C(_06531_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14764_ (.A1(_03457_),
    .A2(_06420_),
    .ZN(_06755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14765_ (.A1(_03458_),
    .A2(_03224_),
    .B(_06755_),
    .ZN(_06756_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14766_ (.A1(_06726_),
    .A2(_06756_),
    .Z(_06757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14767_ (.A1(_06736_),
    .A2(_06752_),
    .ZN(_06758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14768_ (.I(_06741_),
    .Z(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14769_ (.A1(_06735_),
    .A2(_06751_),
    .B(_06759_),
    .ZN(_06760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14770_ (.A1(_06732_),
    .A2(_06758_),
    .B(_06760_),
    .ZN(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14771_ (.A1(_06757_),
    .A2(_06761_),
    .Z(_06762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14772_ (.A1(_06426_),
    .A2(_06762_),
    .ZN(_06763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14773_ (.A1(_03458_),
    .A2(_06532_),
    .B(_06763_),
    .C(_06531_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14774_ (.I(\filters.band[15] ),
    .ZN(_06764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14775_ (.A1(_03470_),
    .A2(_06733_),
    .ZN(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14776_ (.A1(_06764_),
    .A2(_03224_),
    .B(_06765_),
    .ZN(_06766_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14777_ (.A1(_06726_),
    .A2(_06766_),
    .Z(_06767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14778_ (.A1(_06747_),
    .A2(_06756_),
    .ZN(_06768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14779_ (.A1(_06757_),
    .A2(_06761_),
    .ZN(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14780_ (.A1(_06768_),
    .A2(_06769_),
    .ZN(_06770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14781_ (.A1(_06767_),
    .A2(_06770_),
    .Z(_06771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14782_ (.A1(_05570_),
    .A2(_06771_),
    .ZN(_06772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14783_ (.I(_02355_),
    .Z(_06773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _14784_ (.A1(_06764_),
    .A2(_06532_),
    .B(_06772_),
    .C(_06773_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14785_ (.I(_05572_),
    .Z(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14786_ (.A1(_06757_),
    .A2(_06767_),
    .ZN(_06775_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14787_ (.A1(_06758_),
    .A2(_06775_),
    .Z(_06776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14788_ (.A1(_06756_),
    .A2(_06766_),
    .B(_06759_),
    .ZN(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _14789_ (.A1(_06760_),
    .A2(_06775_),
    .B1(_06776_),
    .B2(_06732_),
    .C(_06777_),
    .ZN(_06778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14790_ (.I(_06778_),
    .Z(_06779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14791_ (.I(_06723_),
    .Z(_06780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14792_ (.I(_03474_),
    .Z(_06781_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14793_ (.I0(\filters.low[16] ),
    .I1(\filters.band[16] ),
    .S(_06781_),
    .Z(_06782_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14794_ (.A1(_06780_),
    .A2(_06782_),
    .Z(_06783_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14795_ (.A1(_06779_),
    .A2(_06783_),
    .Z(_06784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14796_ (.A1(_06774_),
    .A2(_06784_),
    .ZN(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14797_ (.I(_04187_),
    .Z(_06786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14798_ (.I(_06786_),
    .Z(_06787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14799_ (.A1(\filters.band[16] ),
    .A2(_06787_),
    .B(_03762_),
    .ZN(_06788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14800_ (.A1(_06785_),
    .A2(_06788_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14801_ (.I(_06741_),
    .Z(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14802_ (.I(_06789_),
    .Z(_06790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14803_ (.I(_06790_),
    .Z(_06791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14804_ (.I(_06791_),
    .Z(_06792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14805_ (.I(_06792_),
    .Z(_06793_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14806_ (.A1(_06793_),
    .A2(_06782_),
    .Z(_06794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14807_ (.A1(_06779_),
    .A2(_06783_),
    .B(_06794_),
    .ZN(_06795_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14808_ (.I0(\filters.low[17] ),
    .I1(\filters.band[17] ),
    .S(_06781_),
    .Z(_06796_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14809_ (.A1(_06780_),
    .A2(_06796_),
    .Z(_06797_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14810_ (.A1(_06795_),
    .A2(_06797_),
    .Z(_06798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14811_ (.A1(\filters.band[17] ),
    .A2(_04188_),
    .B(_06739_),
    .ZN(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14812_ (.A1(_06787_),
    .A2(_06798_),
    .B(_06799_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14813_ (.I(_06712_),
    .Z(_06800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14814_ (.I0(\filters.low[18] ),
    .I1(\filters.band[18] ),
    .S(_06098_),
    .Z(_06801_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14815_ (.A1(_06800_),
    .A2(_06801_),
    .ZN(_06802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _14816_ (.A1(_06782_),
    .A2(_06796_),
    .B(_06789_),
    .ZN(_06803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14817_ (.A1(_06779_),
    .A2(_06783_),
    .A3(_06797_),
    .ZN(_06804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14818_ (.A1(_06803_),
    .A2(_06804_),
    .ZN(_06805_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14819_ (.A1(_06802_),
    .A2(_06805_),
    .ZN(_06806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14820_ (.A1(_06774_),
    .A2(_06806_),
    .ZN(_06807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14821_ (.I(_06786_),
    .Z(_06808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14822_ (.A1(\filters.band[18] ),
    .A2(_06808_),
    .B(_03762_),
    .ZN(_06809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14823_ (.A1(_06807_),
    .A2(_06809_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14824_ (.I0(\filters.low[19] ),
    .I1(\filters.band[19] ),
    .S(_06781_),
    .Z(_06810_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14825_ (.A1(_06729_),
    .A2(_06810_),
    .ZN(_06811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14826_ (.A1(_06803_),
    .A2(_06804_),
    .B(_06802_),
    .ZN(_06812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14827_ (.A1(_06793_),
    .A2(_06801_),
    .B(_06812_),
    .ZN(_06813_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14828_ (.A1(_06811_),
    .A2(_06813_),
    .Z(_06814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14829_ (.A1(_06774_),
    .A2(_06814_),
    .ZN(_06815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14830_ (.A1(\filters.band[19] ),
    .A2(_06808_),
    .B(_03762_),
    .ZN(_06816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14831_ (.A1(_06815_),
    .A2(_06816_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14832_ (.I0(\filters.low[20] ),
    .I1(\filters.band[20] ),
    .S(_03474_),
    .Z(_06817_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14833_ (.A1(_06724_),
    .A2(_06817_),
    .ZN(_06818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14834_ (.A1(_06783_),
    .A2(_06797_),
    .ZN(_06819_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _14835_ (.A1(_06802_),
    .A2(_06819_),
    .A3(_06811_),
    .ZN(_06820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14836_ (.A1(_06801_),
    .A2(_06810_),
    .B(_06759_),
    .ZN(_06821_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _14837_ (.A1(_06802_),
    .A2(_06803_),
    .A3(_06811_),
    .B(_06821_),
    .ZN(_06822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _14838_ (.A1(_06779_),
    .A2(_06820_),
    .B(_06822_),
    .ZN(_06823_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14839_ (.A1(_06818_),
    .A2(_06823_),
    .Z(_06824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14840_ (.A1(_06774_),
    .A2(_06824_),
    .ZN(_06825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14841_ (.I(_03508_),
    .Z(_06826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14842_ (.I(_06826_),
    .Z(_06827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14843_ (.A1(\filters.band[20] ),
    .A2(_06808_),
    .B(_06827_),
    .ZN(_06828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14844_ (.A1(_06825_),
    .A2(_06828_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14845_ (.I(_05572_),
    .Z(_06829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14846_ (.A1(_06818_),
    .A2(_06823_),
    .ZN(_06830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14847_ (.A1(_06793_),
    .A2(_06817_),
    .B(_06830_),
    .ZN(_06831_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14848_ (.I0(\filters.low[21] ),
    .I1(\filters.band[21] ),
    .S(_06098_),
    .Z(_06832_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14849_ (.A1(_06724_),
    .A2(_06832_),
    .ZN(_06833_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14850_ (.A1(_06831_),
    .A2(_06833_),
    .Z(_06834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14851_ (.A1(_06829_),
    .A2(_06834_),
    .ZN(_06835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14852_ (.A1(\filters.band[21] ),
    .A2(_06808_),
    .B(_06827_),
    .ZN(_06836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14853_ (.A1(_06835_),
    .A2(_06836_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14854_ (.I0(\filters.low[22] ),
    .I1(\filters.band[22] ),
    .S(_06098_),
    .Z(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14855_ (.A1(_06800_),
    .A2(_06837_),
    .ZN(_06838_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14856_ (.I(_06838_),
    .ZN(_06839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14857_ (.A1(_06817_),
    .A2(_06832_),
    .B(_06789_),
    .ZN(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _14858_ (.A1(_06818_),
    .A2(_06823_),
    .A3(_06833_),
    .B(_06840_),
    .ZN(_06841_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14859_ (.A1(_06839_),
    .A2(_06841_),
    .Z(_06842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14860_ (.A1(_06829_),
    .A2(_06842_),
    .ZN(_06843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14861_ (.I(_06786_),
    .Z(_06844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14862_ (.A1(\filters.band[22] ),
    .A2(_06844_),
    .B(_06827_),
    .ZN(_06845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14863_ (.A1(_06843_),
    .A2(_06845_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _14864_ (.I(\filters.low[23] ),
    .ZN(_06846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14865_ (.A1(\filters.band[23] ),
    .A2(_06781_),
    .ZN(_06847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14866_ (.A1(_06846_),
    .A2(_03475_),
    .B(_06847_),
    .ZN(_06848_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14867_ (.A1(_06800_),
    .A2(_06848_),
    .ZN(_06849_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14868_ (.A1(_06745_),
    .A2(_06837_),
    .Z(_06850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14869_ (.A1(_06839_),
    .A2(_06841_),
    .B(_06850_),
    .ZN(_06851_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14870_ (.A1(_06849_),
    .A2(_06851_),
    .Z(_06852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14871_ (.A1(_06829_),
    .A2(_06852_),
    .ZN(_06853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14872_ (.A1(\filters.band[23] ),
    .A2(_06844_),
    .B(_06827_),
    .ZN(_06854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14873_ (.A1(_06853_),
    .A2(_06854_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _14874_ (.A1(_06818_),
    .A2(_06833_),
    .A3(_06838_),
    .A4(_06849_),
    .ZN(_06855_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14875_ (.A1(_06820_),
    .A2(_06855_),
    .Z(_06856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14876_ (.A1(_06837_),
    .A2(_06848_),
    .B(_06742_),
    .ZN(_06857_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _14877_ (.A1(_06838_),
    .A2(_06840_),
    .A3(_06849_),
    .B(_06857_),
    .ZN(_06858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _14878_ (.A1(_06822_),
    .A2(_06855_),
    .B1(_06856_),
    .B2(_06778_),
    .C(_06858_),
    .ZN(_06859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14879_ (.I(_06724_),
    .Z(_06860_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _14880_ (.I(\filters.low[24] ),
    .ZN(_06861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14881_ (.A1(\filters.band[24] ),
    .A2(_03476_),
    .ZN(_06862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14882_ (.A1(_06861_),
    .A2(_03476_),
    .B(_06862_),
    .ZN(_06863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14883_ (.A1(_06860_),
    .A2(_06863_),
    .Z(_06864_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14884_ (.A1(_06864_),
    .A2(net31),
    .Z(_06865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14885_ (.A1(\filters.band[24] ),
    .A2(_04188_),
    .B(_06739_),
    .ZN(_06866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14886_ (.A1(_06787_),
    .A2(_06865_),
    .B(_06866_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14887_ (.I(_06864_),
    .ZN(_06867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14888_ (.A1(_06747_),
    .A2(_06863_),
    .ZN(_06868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14889_ (.A1(_06859_),
    .A2(_06867_),
    .B(_06868_),
    .ZN(_06869_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14890_ (.I0(\filters.low[25] ),
    .I1(\filters.band[25] ),
    .S(_03475_),
    .Z(_06870_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14891_ (.A1(_06860_),
    .A2(_06870_),
    .Z(_06871_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14892_ (.A1(_06869_),
    .A2(_06871_),
    .Z(_06872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14893_ (.A1(_06829_),
    .A2(_06872_),
    .ZN(_06873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14894_ (.I(_06826_),
    .Z(_06874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14895_ (.A1(\filters.band[25] ),
    .A2(_06844_),
    .B(_06874_),
    .ZN(_06875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14896_ (.A1(_06873_),
    .A2(_06875_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14897_ (.I(_05572_),
    .Z(_06876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14898_ (.I(_06729_),
    .Z(_06877_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14899_ (.I0(\filters.low[26] ),
    .I1(_06495_),
    .S(_03475_),
    .Z(_06878_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14900_ (.A1(_06877_),
    .A2(_06878_),
    .Z(_06879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14901_ (.A1(_06864_),
    .A2(_06871_),
    .ZN(_06880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14902_ (.A1(_06863_),
    .A2(_06870_),
    .B(_06743_),
    .ZN(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14903_ (.A1(_06859_),
    .A2(_06880_),
    .B(_06881_),
    .ZN(_06882_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14904_ (.A1(_06879_),
    .A2(_06882_),
    .Z(_06883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14905_ (.A1(_06876_),
    .A2(_06883_),
    .ZN(_06884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14906_ (.A1(_06495_),
    .A2(_06844_),
    .B(_06874_),
    .ZN(_06885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14907_ (.A1(_06884_),
    .A2(_06885_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14908_ (.I(_06729_),
    .Z(_06886_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14909_ (.I0(\filters.low[27] ),
    .I1(_06544_),
    .S(_03476_),
    .Z(_06887_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14910_ (.A1(_06886_),
    .A2(_06887_),
    .Z(_06888_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14911_ (.A1(_06792_),
    .A2(_06878_),
    .Z(_06889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14912_ (.A1(_06879_),
    .A2(_06882_),
    .B(_06889_),
    .ZN(_06890_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14913_ (.A1(_06888_),
    .A2(_06890_),
    .ZN(_06891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14914_ (.A1(_06876_),
    .A2(_06891_),
    .ZN(_06892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14915_ (.I(_06786_),
    .Z(_06893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14916_ (.A1(_06544_),
    .A2(_06893_),
    .B(_06874_),
    .ZN(_06894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14917_ (.A1(_06892_),
    .A2(_06894_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14918_ (.A1(_06879_),
    .A2(_06888_),
    .ZN(_06895_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _14919_ (.A1(_06880_),
    .A2(_06895_),
    .Z(_06896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14920_ (.A1(_06878_),
    .A2(_06887_),
    .B(_06743_),
    .ZN(_06897_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _14921_ (.A1(_06881_),
    .A2(_06895_),
    .B1(_06896_),
    .B2(_06859_),
    .C(_06897_),
    .ZN(_06898_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _14922_ (.I(\filters.low[28] ),
    .ZN(_06899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14923_ (.A1(_06639_),
    .A2(_03477_),
    .ZN(_06900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14924_ (.A1(_06899_),
    .A2(_03478_),
    .B(_06900_),
    .ZN(_06901_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14925_ (.A1(_06790_),
    .A2(_06901_),
    .Z(_06902_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14926_ (.A1(_06898_),
    .A2(_06902_),
    .Z(_06903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14927_ (.A1(_06876_),
    .A2(_06903_),
    .ZN(_06904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14928_ (.A1(_06639_),
    .A2(_06893_),
    .B(_06874_),
    .ZN(_06905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14929_ (.A1(_06904_),
    .A2(_06905_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _14930_ (.I(\filters.low[29] ),
    .ZN(_06906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14931_ (.A1(_06568_),
    .A2(_03477_),
    .ZN(_06907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _14932_ (.A1(_06906_),
    .A2(_03477_),
    .B(_06907_),
    .ZN(_06908_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _14933_ (.A1(_06743_),
    .A2(_06908_),
    .ZN(_06909_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14934_ (.A1(_06744_),
    .A2(_06901_),
    .Z(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14935_ (.A1(_06898_),
    .A2(_06902_),
    .B(_06910_),
    .ZN(_06911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14936_ (.A1(_06909_),
    .A2(_06911_),
    .Z(_06912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14937_ (.A1(_06876_),
    .A2(_06912_),
    .ZN(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14938_ (.I(_06826_),
    .Z(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14939_ (.A1(_06568_),
    .A2(_06893_),
    .B(_06914_),
    .ZN(_06915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14940_ (.A1(_06913_),
    .A2(_06915_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _14941_ (.I(\filters.low[30] ),
    .ZN(_06916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14942_ (.A1(\filters.band[30] ),
    .A2(_03478_),
    .ZN(_06917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14943_ (.A1(_06916_),
    .A2(_03479_),
    .B(_06917_),
    .ZN(_06918_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14944_ (.I(_06902_),
    .ZN(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14945_ (.A1(_06919_),
    .A2(_06909_),
    .ZN(_06920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _14946_ (.A1(_06792_),
    .A2(_06908_),
    .B1(_06920_),
    .B2(_06898_),
    .C(_06910_),
    .ZN(_06921_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14947_ (.A1(_06747_),
    .A2(_06918_),
    .A3(_06921_),
    .ZN(_06922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14948_ (.A1(_05573_),
    .A2(_06922_),
    .ZN(_06923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14949_ (.A1(\filters.band[30] ),
    .A2(_06893_),
    .B(_06914_),
    .ZN(_06924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14950_ (.A1(_06923_),
    .A2(_06924_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14951_ (.A1(_06745_),
    .A2(_06918_),
    .ZN(_06925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14952_ (.A1(_06745_),
    .A2(_06918_),
    .ZN(_06926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14953_ (.A1(_06925_),
    .A2(_06921_),
    .B(_06926_),
    .ZN(_06927_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14954_ (.I0(\filters.low[31] ),
    .I1(\filters.band[31] ),
    .S(_03479_),
    .Z(_06928_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14955_ (.A1(_06793_),
    .A2(_06927_),
    .A3(_06928_),
    .ZN(_06929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14956_ (.A1(\filters.band[31] ),
    .A2(_04188_),
    .B(_06739_),
    .ZN(_06930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14957_ (.A1(_06787_),
    .A2(_06929_),
    .B(_06930_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14958_ (.A1(_03758_),
    .A2(_04198_),
    .ZN(_06931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14959_ (.I(_06931_),
    .Z(_06932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14960_ (.I(_06932_),
    .Z(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14961_ (.I(_06933_),
    .Z(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14962_ (.I(\filters.low[0] ),
    .ZN(_06935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14963_ (.A1(_04583_),
    .A2(_04720_),
    .Z(_06936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14964_ (.I(_06932_),
    .Z(_06937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14965_ (.A1(_06935_),
    .A2(_06936_),
    .B(_06937_),
    .ZN(_06938_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _14966_ (.A1(_04583_),
    .A2(_04720_),
    .ZN(_06939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14967_ (.A1(_05561_),
    .A2(_06939_),
    .ZN(_06940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14968_ (.I(_03561_),
    .Z(_06941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _14969_ (.A1(_04243_),
    .A2(_06934_),
    .B1(_06938_),
    .B2(_06940_),
    .C(_06941_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14970_ (.I(_01944_),
    .Z(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14971_ (.I(_06932_),
    .Z(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14972_ (.A1(_04583_),
    .A2(_04720_),
    .B(_04721_),
    .ZN(_06944_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _14973_ (.A1(_04458_),
    .A2(_04545_),
    .A3(_06944_),
    .ZN(_06945_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _14974_ (.A1(_01769_),
    .A2(_01755_),
    .A3(\channels.sample1[0] ),
    .A4(\channels.sample2[0] ),
    .Z(_06946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _14975_ (.A1(_01755_),
    .A2(\channels.sample1[0] ),
    .B1(\channels.sample2[0] ),
    .B2(_01769_),
    .ZN(_06947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14976_ (.A1(_06946_),
    .A2(_06947_),
    .ZN(_06948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14977_ (.A1(_01778_),
    .A2(\channels.sample3[0] ),
    .ZN(_06949_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _14978_ (.A1(_05676_),
    .A2(_06948_),
    .A3(_06949_),
    .ZN(_06950_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14979_ (.I(_06950_),
    .ZN(_06951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14980_ (.A1(_06935_),
    .A2(_06936_),
    .B(_06951_),
    .ZN(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14981_ (.A1(_05561_),
    .A2(_06939_),
    .A3(_06950_),
    .ZN(_06953_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14982_ (.A1(_06945_),
    .A2(_06952_),
    .A3(_06953_),
    .ZN(_06954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14983_ (.A1(_06952_),
    .A2(_06953_),
    .B(_06945_),
    .ZN(_06955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14984_ (.A1(_06933_),
    .A2(_06955_),
    .ZN(_06956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14985_ (.A1(\filters.high[1] ),
    .A2(_06943_),
    .B1(_06954_),
    .B2(_06956_),
    .ZN(_06957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14986_ (.A1(_06942_),
    .A2(_06957_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _14987_ (.I(_06932_),
    .Z(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _14988_ (.A1(_06952_),
    .A2(_06954_),
    .Z(_06959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14989_ (.A1(_06946_),
    .A2(_06947_),
    .B(_06949_),
    .ZN(_06960_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14990_ (.A1(_01783_),
    .A2(\channels.sample3[0] ),
    .A3(_06948_),
    .ZN(_06961_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _14991_ (.A1(_05676_),
    .A2(_06960_),
    .A3(_06961_),
    .ZN(_06962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14992_ (.A1(_04546_),
    .A2(_04722_),
    .ZN(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _14993_ (.A1(_01768_),
    .A2(_01754_),
    .A3(\channels.sample1[1] ),
    .A4(\channels.sample2[1] ),
    .Z(_06964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14994_ (.A1(_01754_),
    .A2(\channels.sample1[1] ),
    .B1(\channels.sample2[1] ),
    .B2(_01768_),
    .ZN(_06965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14995_ (.A1(_06964_),
    .A2(_06965_),
    .ZN(_06966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14996_ (.A1(_01778_),
    .A2(\channels.sample3[1] ),
    .ZN(_06967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14997_ (.A1(_06966_),
    .A2(_06967_),
    .Z(_06968_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _14998_ (.A1(_06946_),
    .A2(_06947_),
    .A3(_06949_),
    .ZN(_06969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14999_ (.A1(_06946_),
    .A2(_06969_),
    .ZN(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15000_ (.A1(_06968_),
    .A2(_06970_),
    .Z(_06971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15001_ (.A1(\filters.low[2] ),
    .A2(_06971_),
    .Z(_06972_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15002_ (.A1(_06963_),
    .A2(_05061_),
    .A3(_06972_),
    .Z(_06973_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _15003_ (.A1(_06962_),
    .A2(_06973_),
    .ZN(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15004_ (.A1(_06959_),
    .A2(_06974_),
    .Z(_06975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15005_ (.I(_06931_),
    .Z(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15006_ (.A1(_06959_),
    .A2(_06974_),
    .B(_06976_),
    .ZN(_06977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15007_ (.A1(\filters.high[2] ),
    .A2(_06958_),
    .B1(_06975_),
    .B2(_06977_),
    .ZN(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15008_ (.A1(_06942_),
    .A2(_06978_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15009_ (.I(_06976_),
    .Z(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15010_ (.A1(\filters.high[3] ),
    .A2(_06979_),
    .ZN(_06980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15011_ (.A1(_06962_),
    .A2(_06973_),
    .ZN(_06981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _15012_ (.A1(_06959_),
    .A2(_06974_),
    .B(_06981_),
    .ZN(_06982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15013_ (.A1(_06968_),
    .A2(_06970_),
    .ZN(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15014_ (.I(_06967_),
    .ZN(_06984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15015_ (.A1(_06966_),
    .A2(_06984_),
    .B(_06964_),
    .ZN(_06985_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _15016_ (.A1(\filters.filt_2 ),
    .A2(\filters.filt_1 ),
    .A3(\channels.sample1[2] ),
    .A4(\channels.sample2[2] ),
    .Z(_06986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15017_ (.A1(\filters.filt_1 ),
    .A2(\channels.sample1[2] ),
    .B1(\channels.sample2[2] ),
    .B2(\filters.filt_2 ),
    .ZN(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15018_ (.A1(_06986_),
    .A2(_06987_),
    .Z(_06988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15019_ (.A1(\filters.filt_3 ),
    .A2(\channels.sample3[2] ),
    .ZN(_06989_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15020_ (.A1(_06988_),
    .A2(_06989_),
    .ZN(_06990_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15021_ (.A1(_06985_),
    .A2(_06990_),
    .ZN(_06991_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15022_ (.A1(_06983_),
    .A2(_06991_),
    .ZN(_06992_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15023_ (.A1(\filters.low[3] ),
    .A2(_06992_),
    .Z(_06993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15024_ (.A1(_06963_),
    .A2(_05061_),
    .B(_05066_),
    .ZN(_06994_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15025_ (.A1(net38),
    .A2(_06993_),
    .A3(_06994_),
    .Z(_06995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15026_ (.A1(_06963_),
    .A2(_05061_),
    .Z(_06996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15027_ (.A1(_03270_),
    .A2(_06971_),
    .ZN(_06997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15028_ (.A1(_06972_),
    .A2(_06996_),
    .B(_06997_),
    .ZN(_06998_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15029_ (.A1(_06995_),
    .A2(_06998_),
    .Z(_06999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15030_ (.A1(_06982_),
    .A2(_06999_),
    .B(_06976_),
    .ZN(_07000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15031_ (.A1(_06982_),
    .A2(_06999_),
    .B(_07000_),
    .ZN(_07001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15032_ (.A1(_06980_),
    .A2(_07001_),
    .B(_03750_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15033_ (.A1(\filters.high[4] ),
    .A2(_06979_),
    .ZN(_07002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15034_ (.A1(_03497_),
    .A2(_04809_),
    .ZN(_07003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15035_ (.I(_07003_),
    .Z(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15036_ (.I(_07004_),
    .Z(_07005_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _15037_ (.A1(_06968_),
    .A2(_06970_),
    .A3(_06991_),
    .B1(_06990_),
    .B2(_06985_),
    .ZN(_07006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15038_ (.A1(_06988_),
    .A2(_06989_),
    .ZN(_07007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15039_ (.A1(_06986_),
    .A2(_07007_),
    .ZN(_07008_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _15040_ (.A1(\filters.filt_2 ),
    .A2(\filters.filt_1 ),
    .A3(\channels.sample1[3] ),
    .A4(\channels.sample2[3] ),
    .Z(_07009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15041_ (.A1(_01754_),
    .A2(\channels.sample1[3] ),
    .B1(\channels.sample2[3] ),
    .B2(_01768_),
    .ZN(_07010_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15042_ (.A1(_07009_),
    .A2(_07010_),
    .Z(_07011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15043_ (.A1(_01778_),
    .A2(\channels.sample3[3] ),
    .ZN(_07012_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15044_ (.A1(_07011_),
    .A2(_07012_),
    .ZN(_07013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15045_ (.A1(_07008_),
    .A2(_07013_),
    .Z(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15046_ (.A1(_07006_),
    .A2(_07014_),
    .Z(_07015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15047_ (.I(_05042_),
    .ZN(_07016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15048_ (.A1(_04723_),
    .A2(_05062_),
    .B(_05068_),
    .ZN(_07017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15049_ (.A1(_07016_),
    .A2(_07017_),
    .Z(_07018_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _15050_ (.A1(\filters.low[4] ),
    .A2(_07015_),
    .A3(_07018_),
    .ZN(_07019_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15051_ (.A1(net38),
    .A2(_06994_),
    .ZN(_07020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15052_ (.A1(_03284_),
    .A2(_06992_),
    .ZN(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15053_ (.A1(_06993_),
    .A2(_07020_),
    .B(_07021_),
    .ZN(_07022_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _15054_ (.A1(_07019_),
    .A2(_07022_),
    .ZN(_07023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15055_ (.A1(_06995_),
    .A2(_06998_),
    .ZN(_07024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _15056_ (.A1(_06982_),
    .A2(_06999_),
    .B(_07024_),
    .ZN(_07025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15057_ (.A1(_07023_),
    .A2(_07025_),
    .Z(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15058_ (.A1(_07005_),
    .A2(_07026_),
    .ZN(_07027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15059_ (.A1(_07002_),
    .A2(_07027_),
    .B(_03750_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15060_ (.A1(_07019_),
    .A2(_07022_),
    .Z(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15061_ (.A1(_07023_),
    .A2(_07025_),
    .B(_07028_),
    .ZN(_07029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15062_ (.A1(_05994_),
    .A2(_07015_),
    .ZN(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15063_ (.A1(_05994_),
    .A2(_07015_),
    .ZN(_07031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15064_ (.A1(_07030_),
    .A2(_07018_),
    .B(_07031_),
    .ZN(_07032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15065_ (.A1(_05040_),
    .A2(_05072_),
    .B(_05019_),
    .ZN(_07033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15066_ (.A1(_07016_),
    .A2(_07017_),
    .B(_07033_),
    .ZN(_07034_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15067_ (.A1(_07008_),
    .A2(_07013_),
    .Z(_07035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15068_ (.A1(_07006_),
    .A2(_07014_),
    .ZN(_07036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15069_ (.A1(_07035_),
    .A2(_07036_),
    .Z(_07037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15070_ (.A1(_07011_),
    .A2(_07012_),
    .ZN(_07038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15071_ (.A1(_07009_),
    .A2(_07038_),
    .ZN(_07039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15072_ (.A1(_01779_),
    .A2(\channels.sample3[4] ),
    .ZN(_07040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15073_ (.A1(_01770_),
    .A2(\channels.sample2[4] ),
    .ZN(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15074_ (.A1(_01756_),
    .A2(\channels.sample1[4] ),
    .ZN(_07042_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15075_ (.A1(_07040_),
    .A2(_07041_),
    .A3(_07042_),
    .Z(_07043_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _15076_ (.A1(_07037_),
    .A2(_07039_),
    .A3(_07043_),
    .ZN(_07044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15077_ (.A1(\filters.low[5] ),
    .A2(_07044_),
    .Z(_07045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15078_ (.I(_07045_),
    .ZN(_07046_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15079_ (.A1(_05018_),
    .A2(_07034_),
    .A3(_07046_),
    .Z(_07047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15080_ (.A1(_07032_),
    .A2(_07047_),
    .ZN(_07048_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15081_ (.A1(_07032_),
    .A2(_07047_),
    .Z(_07049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15082_ (.A1(_07048_),
    .A2(_07049_),
    .ZN(_07050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15083_ (.I(_07003_),
    .Z(_07051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15084_ (.I(_07051_),
    .Z(_07052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15085_ (.A1(_07029_),
    .A2(_07050_),
    .B(_07052_),
    .ZN(_07053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15086_ (.A1(_07029_),
    .A2(_07050_),
    .B(_07053_),
    .ZN(_07054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15087_ (.I(_07051_),
    .Z(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15088_ (.A1(\filters.high[5] ),
    .A2(_07055_),
    .B(_06914_),
    .ZN(_07056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15089_ (.A1(_07054_),
    .A2(_07056_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15090_ (.I(_07051_),
    .Z(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15091_ (.I(_07057_),
    .Z(_07058_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _15092_ (.A1(_07023_),
    .A2(_07025_),
    .B(_07049_),
    .C(_07028_),
    .ZN(_07059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15093_ (.A1(_07048_),
    .A2(_07059_),
    .ZN(_07060_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15094_ (.A1(_07039_),
    .A2(_07043_),
    .Z(_07061_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15095_ (.A1(_07039_),
    .A2(_07043_),
    .Z(_07062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15096_ (.A1(_07037_),
    .A2(_07061_),
    .B(_07062_),
    .ZN(_07063_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15097_ (.A1(_07041_),
    .A2(_07042_),
    .Z(_07064_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15098_ (.A1(_07041_),
    .A2(_07042_),
    .Z(_07065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15099_ (.A1(_07040_),
    .A2(_07064_),
    .B(_07065_),
    .ZN(_07066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15100_ (.A1(_01779_),
    .A2(\channels.sample3[5] ),
    .ZN(_07067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15101_ (.A1(_01769_),
    .A2(\channels.sample2[5] ),
    .ZN(_07068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15102_ (.A1(_01755_),
    .A2(\channels.sample1[5] ),
    .ZN(_07069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15103_ (.A1(_07068_),
    .A2(_07069_),
    .Z(_07070_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15104_ (.A1(_07067_),
    .A2(_07070_),
    .Z(_07071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15105_ (.I(_07071_),
    .ZN(_07072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15106_ (.A1(_07066_),
    .A2(_07072_),
    .Z(_07073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15107_ (.A1(_07063_),
    .A2(_07073_),
    .Z(_07074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15108_ (.A1(\filters.low[6] ),
    .A2(_07074_),
    .Z(_07075_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _15109_ (.A1(net65),
    .A2(_05069_),
    .A3(_05074_),
    .ZN(_07076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15110_ (.A1(_07076_),
    .A2(_05450_),
    .Z(_07077_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15111_ (.A1(_07075_),
    .A2(_07077_),
    .Z(_07078_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15112_ (.A1(_05018_),
    .A2(_07034_),
    .ZN(_07079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15113_ (.A1(_03312_),
    .A2(_07044_),
    .ZN(_07080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15114_ (.I(_07080_),
    .ZN(_07081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15115_ (.A1(_07079_),
    .A2(_07046_),
    .B(_07081_),
    .ZN(_07082_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15116_ (.A1(_07078_),
    .A2(_07082_),
    .Z(_07083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15117_ (.A1(_07060_),
    .A2(_07083_),
    .Z(_07084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15118_ (.I(_07004_),
    .Z(_07085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15119_ (.I(_06738_),
    .Z(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15120_ (.A1(\filters.high[6] ),
    .A2(_07085_),
    .B(_07086_),
    .ZN(_07087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15121_ (.A1(_07058_),
    .A2(_07084_),
    .B(_07087_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15122_ (.I(_06937_),
    .Z(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15123_ (.A1(_05446_),
    .A2(_05449_),
    .Z(_07089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15124_ (.A1(_07076_),
    .A2(_05450_),
    .B(_07089_),
    .ZN(_07090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15125_ (.A1(_07066_),
    .A2(_07072_),
    .ZN(_07091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15126_ (.A1(_07063_),
    .A2(_07073_),
    .ZN(_07092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15127_ (.A1(_07091_),
    .A2(_07092_),
    .ZN(_07093_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15128_ (.A1(_01780_),
    .A2(_01939_),
    .A3(_07070_),
    .ZN(_07094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15129_ (.A1(_07068_),
    .A2(_07069_),
    .B(_07094_),
    .ZN(_07095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15130_ (.I(_07095_),
    .ZN(_07096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15131_ (.A1(_01779_),
    .A2(\channels.sample3[6] ),
    .ZN(_07097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15132_ (.A1(_01770_),
    .A2(\channels.sample2[6] ),
    .ZN(_07098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15133_ (.A1(_01756_),
    .A2(\channels.sample1[6] ),
    .ZN(_07099_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15134_ (.A1(_07097_),
    .A2(_07098_),
    .A3(_07099_),
    .Z(_07100_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15135_ (.A1(_07093_),
    .A2(_07096_),
    .A3(_07100_),
    .Z(_07101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15136_ (.A1(\filters.low[7] ),
    .A2(_07101_),
    .Z(_07102_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15137_ (.A1(_05445_),
    .A2(_07090_),
    .A3(_07102_),
    .Z(_07103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15138_ (.A1(_03331_),
    .A2(_07074_),
    .ZN(_07104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15139_ (.A1(_07075_),
    .A2(_07077_),
    .B(_07104_),
    .ZN(_07105_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15140_ (.A1(_07103_),
    .A2(_07105_),
    .Z(_07106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15141_ (.A1(_07078_),
    .A2(_07082_),
    .ZN(_07107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15142_ (.A1(_07048_),
    .A2(_07059_),
    .A3(_07083_),
    .ZN(_07108_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15143_ (.A1(_07107_),
    .A2(_07108_),
    .Z(_07109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15144_ (.I(_07051_),
    .Z(_07110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15145_ (.A1(_07106_),
    .A2(_07109_),
    .B(_07110_),
    .ZN(_07111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15146_ (.A1(_07106_),
    .A2(_07109_),
    .B(_07111_),
    .ZN(_07112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15147_ (.A1(_03345_),
    .A2(_07088_),
    .B(_07112_),
    .C(_06773_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15148_ (.A1(_07078_),
    .A2(_07082_),
    .Z(_07113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15149_ (.A1(_07103_),
    .A2(_07105_),
    .ZN(_07114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15150_ (.A1(_07103_),
    .A2(_07105_),
    .ZN(_07115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15151_ (.A1(_07113_),
    .A2(_07114_),
    .B(_07115_),
    .ZN(_07116_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _15152_ (.A1(_07048_),
    .A2(_07059_),
    .A3(_07083_),
    .A4(_07106_),
    .ZN(_07117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15153_ (.A1(_07116_),
    .A2(_07117_),
    .ZN(_07118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15154_ (.A1(_05456_),
    .A2(_05457_),
    .ZN(_07119_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _15155_ (.A1(_07076_),
    .A2(_05445_),
    .A3(_05450_),
    .B(_07119_),
    .ZN(_07120_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15156_ (.A1(_05433_),
    .A2(_07120_),
    .ZN(_07121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15157_ (.A1(_07096_),
    .A2(_07100_),
    .ZN(_07122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15158_ (.A1(_07096_),
    .A2(_07100_),
    .ZN(_07123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15159_ (.A1(_07093_),
    .A2(_07122_),
    .B(_07123_),
    .ZN(_07124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15160_ (.I(_07097_),
    .ZN(_07125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15161_ (.A1(_07098_),
    .A2(_07099_),
    .ZN(_07126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15162_ (.A1(_07098_),
    .A2(_07099_),
    .ZN(_07127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15163_ (.A1(_07125_),
    .A2(_07126_),
    .B(_07127_),
    .ZN(_07128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15164_ (.A1(_01780_),
    .A2(\channels.sample3[7] ),
    .ZN(_07129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15165_ (.A1(_01770_),
    .A2(\channels.sample2[7] ),
    .ZN(_07130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15166_ (.A1(_01756_),
    .A2(\channels.sample1[7] ),
    .ZN(_07131_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15167_ (.A1(_07130_),
    .A2(_07131_),
    .Z(_07132_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15168_ (.A1(_07129_),
    .A2(_07132_),
    .Z(_07133_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _15169_ (.A1(_07124_),
    .A2(_07128_),
    .A3(_07133_),
    .ZN(_07134_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15170_ (.A1(\filters.low[8] ),
    .A2(_07134_),
    .ZN(_07135_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15171_ (.A1(_07121_),
    .A2(_07135_),
    .Z(_07136_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15172_ (.A1(_05445_),
    .A2(_07090_),
    .ZN(_07137_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15173_ (.A1(_03347_),
    .A2(_07101_),
    .Z(_07138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15174_ (.I(_07138_),
    .ZN(_07139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _15175_ (.A1(_07137_),
    .A2(_07102_),
    .B(_07139_),
    .ZN(_07140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15176_ (.A1(_07136_),
    .A2(_07140_),
    .Z(_07141_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15177_ (.A1(_07118_),
    .A2(_07141_),
    .Z(_07142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15178_ (.A1(_06937_),
    .A2(_07142_),
    .ZN(_07143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15179_ (.A1(_03361_),
    .A2(_07088_),
    .B(_07143_),
    .C(_06773_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15180_ (.A1(_05408_),
    .A2(_05432_),
    .ZN(_07144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15181_ (.A1(_07144_),
    .A2(_07120_),
    .B(_05454_),
    .ZN(_07145_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15182_ (.A1(_07128_),
    .A2(_07133_),
    .Z(_07146_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15183_ (.A1(_07128_),
    .A2(_07133_),
    .Z(_07147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15184_ (.A1(_07124_),
    .A2(_07146_),
    .B(_07147_),
    .ZN(_07148_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15185_ (.A1(_01781_),
    .A2(_01989_),
    .A3(_07132_),
    .ZN(_07149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15186_ (.A1(_07130_),
    .A2(_07131_),
    .B(_07149_),
    .ZN(_07150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15187_ (.I(_07150_),
    .ZN(_07151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15188_ (.A1(_01780_),
    .A2(\channels.sample3[8] ),
    .ZN(_07152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15189_ (.A1(_01771_),
    .A2(\channels.sample2[8] ),
    .ZN(_07153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15190_ (.A1(_01757_),
    .A2(\channels.sample1[8] ),
    .ZN(_07154_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15191_ (.A1(_07152_),
    .A2(_07153_),
    .A3(_07154_),
    .Z(_07155_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15192_ (.A1(_07148_),
    .A2(_07151_),
    .A3(_07155_),
    .Z(_07156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15193_ (.A1(\filters.low[9] ),
    .A2(_07156_),
    .ZN(_07157_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _15194_ (.A1(_05407_),
    .A2(_07145_),
    .A3(_07157_),
    .Z(_07158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15195_ (.I(_07135_),
    .ZN(_07159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15196_ (.A1(_03362_),
    .A2(_07134_),
    .ZN(_07160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15197_ (.A1(_07121_),
    .A2(_07159_),
    .B(_07160_),
    .ZN(_07161_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15198_ (.A1(_07158_),
    .A2(_07161_),
    .Z(_07162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15199_ (.A1(_07136_),
    .A2(_07140_),
    .ZN(_07163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15200_ (.A1(_07118_),
    .A2(_07141_),
    .B(_07163_),
    .ZN(_07164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15201_ (.A1(_07162_),
    .A2(_07164_),
    .B(_07110_),
    .ZN(_07165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15202_ (.A1(_07162_),
    .A2(_07164_),
    .B(_07165_),
    .ZN(_07166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15203_ (.A1(_03375_),
    .A2(_07088_),
    .B(_07166_),
    .C(_06773_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15204_ (.A1(_07136_),
    .A2(_07140_),
    .ZN(_07167_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15205_ (.A1(_07161_),
    .A2(_07158_),
    .ZN(_07168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _15206_ (.A1(_07116_),
    .A2(_07117_),
    .B(_07167_),
    .C(_07168_),
    .ZN(_07169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15207_ (.A1(_07158_),
    .A2(_07161_),
    .ZN(_07170_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _15208_ (.A1(_07136_),
    .A2(_07140_),
    .B1(_07158_),
    .B2(_07161_),
    .ZN(_07171_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _15209_ (.A1(_07170_),
    .A2(_07171_),
    .Z(_07172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15210_ (.A1(_07151_),
    .A2(_07155_),
    .ZN(_07173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15211_ (.A1(_07151_),
    .A2(_07155_),
    .ZN(_07174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15212_ (.A1(_07148_),
    .A2(_07173_),
    .B(_07174_),
    .ZN(_07175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15213_ (.I(_07152_),
    .ZN(_07176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15214_ (.A1(_07153_),
    .A2(_07154_),
    .ZN(_07177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15215_ (.A1(_07153_),
    .A2(_07154_),
    .ZN(_07178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15216_ (.A1(_07176_),
    .A2(_07177_),
    .B(_07178_),
    .ZN(_07179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15217_ (.A1(_01781_),
    .A2(\channels.sample3[9] ),
    .ZN(_07180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15218_ (.A1(_01771_),
    .A2(\channels.sample2[9] ),
    .ZN(_07181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15219_ (.A1(_01757_),
    .A2(\channels.sample1[9] ),
    .ZN(_07182_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15220_ (.A1(_07181_),
    .A2(_07182_),
    .Z(_07183_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15221_ (.A1(_07180_),
    .A2(_07183_),
    .Z(_07184_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _15222_ (.A1(_07175_),
    .A2(_07179_),
    .A3(_07184_),
    .ZN(_07185_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15223_ (.A1(\filters.low[10] ),
    .A2(_05559_),
    .A3(_07185_),
    .Z(_07186_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15224_ (.I(_07186_),
    .ZN(_07187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15225_ (.A1(_05407_),
    .A2(_07145_),
    .Z(_07188_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15226_ (.I(_07157_),
    .ZN(_07189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15227_ (.A1(_03376_),
    .A2(_07156_),
    .ZN(_07190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _15228_ (.A1(_07188_),
    .A2(_07189_),
    .B(_07190_),
    .ZN(_07191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15229_ (.A1(_07187_),
    .A2(_07191_),
    .Z(_07192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15230_ (.A1(_07169_),
    .A2(_07172_),
    .B(_07192_),
    .ZN(_07193_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _15231_ (.A1(_07192_),
    .A2(_07169_),
    .A3(_07172_),
    .ZN(_07194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15232_ (.A1(_06933_),
    .A2(_07194_),
    .ZN(_07195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15233_ (.A1(\filters.high[10] ),
    .A2(_06958_),
    .B1(_07193_),
    .B2(_07195_),
    .ZN(_07196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15234_ (.A1(_06942_),
    .A2(_07196_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15235_ (.A1(_03396_),
    .A2(_07185_),
    .ZN(_07197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15236_ (.A1(_03396_),
    .A2(_07185_),
    .ZN(_07198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15237_ (.A1(_05560_),
    .A2(_07197_),
    .B(_07198_),
    .ZN(_07199_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15238_ (.A1(_07179_),
    .A2(_07184_),
    .Z(_07200_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15239_ (.A1(_07179_),
    .A2(_07184_),
    .Z(_07201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15240_ (.A1(_07175_),
    .A2(_07200_),
    .B(_07201_),
    .ZN(_07202_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15241_ (.A1(_01782_),
    .A2(_02040_),
    .A3(_07183_),
    .ZN(_07203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15242_ (.A1(_07181_),
    .A2(_07182_),
    .B(_07203_),
    .ZN(_07204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15243_ (.I(_07204_),
    .ZN(_07205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15244_ (.A1(_01781_),
    .A2(\channels.sample3[10] ),
    .ZN(_07206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15245_ (.A1(_01772_),
    .A2(\channels.sample2[10] ),
    .ZN(_07207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15246_ (.A1(_01758_),
    .A2(\channels.sample1[10] ),
    .ZN(_07208_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15247_ (.A1(_07206_),
    .A2(_07207_),
    .A3(_07208_),
    .Z(_07209_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15248_ (.A1(_07202_),
    .A2(_07205_),
    .A3(_07209_),
    .Z(_07210_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15249_ (.A1(\filters.low[11] ),
    .A2(_07210_),
    .Z(_07211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15250_ (.A1(_03413_),
    .A2(_07210_),
    .ZN(_07212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15251_ (.A1(_07211_),
    .A2(_07212_),
    .ZN(_07213_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _15252_ (.A1(_07213_),
    .A2(_05675_),
    .ZN(_07214_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15253_ (.A1(_07199_),
    .A2(_07214_),
    .ZN(_07215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15254_ (.A1(_07187_),
    .A2(_07191_),
    .B(_07193_),
    .ZN(_07216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15255_ (.A1(_07215_),
    .A2(_07216_),
    .B(_07110_),
    .ZN(_07217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15256_ (.A1(_07215_),
    .A2(_07216_),
    .B(_07217_),
    .ZN(_07218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15257_ (.I(_02355_),
    .Z(_07219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15258_ (.A1(_03412_),
    .A2(_07088_),
    .B(_07218_),
    .C(_07219_),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15259_ (.A1(_07199_),
    .A2(_07214_),
    .Z(_07220_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15260_ (.A1(_07169_),
    .A2(_07172_),
    .B(_07220_),
    .C(_07192_),
    .ZN(_07221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15261_ (.A1(_07187_),
    .A2(_07191_),
    .ZN(_07222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15262_ (.A1(_07199_),
    .A2(_07214_),
    .ZN(_07223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15263_ (.A1(_07199_),
    .A2(_07214_),
    .ZN(_07224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15264_ (.A1(_07222_),
    .A2(_07223_),
    .B(_07224_),
    .ZN(_07225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15265_ (.A1(_07221_),
    .A2(_07225_),
    .ZN(_07226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15266_ (.I(_07226_),
    .ZN(_07227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15267_ (.A1(_07205_),
    .A2(_07209_),
    .ZN(_07228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15268_ (.A1(_07205_),
    .A2(_07209_),
    .ZN(_07229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15269_ (.A1(_07202_),
    .A2(_07228_),
    .B(_07229_),
    .ZN(_07230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15270_ (.I(_07206_),
    .ZN(_07231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15271_ (.A1(_07207_),
    .A2(_07208_),
    .ZN(_07232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15272_ (.A1(_07207_),
    .A2(_07208_),
    .ZN(_07233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15273_ (.A1(_07231_),
    .A2(_07232_),
    .B(_07233_),
    .ZN(_07234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15274_ (.A1(_01782_),
    .A2(\channels.sample3[11] ),
    .ZN(_07235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15275_ (.A1(_01771_),
    .A2(\channels.sample2[11] ),
    .ZN(_07236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15276_ (.A1(_01757_),
    .A2(\channels.sample1[11] ),
    .ZN(_07237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15277_ (.A1(_07236_),
    .A2(_07237_),
    .Z(_07238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15278_ (.A1(_07235_),
    .A2(_07238_),
    .Z(_07239_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _15279_ (.A1(_07230_),
    .A2(_07234_),
    .A3(_07239_),
    .ZN(_07240_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15280_ (.A1(\filters.low[12] ),
    .A2(_07240_),
    .Z(_07241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15281_ (.A1(_03424_),
    .A2(_07240_),
    .ZN(_07242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15282_ (.A1(_07241_),
    .A2(_07242_),
    .ZN(_07243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15283_ (.A1(_05675_),
    .A2(_07213_),
    .B(_07211_),
    .ZN(_07244_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15284_ (.A1(_05779_),
    .A2(_07243_),
    .A3(_07244_),
    .Z(_07245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15285_ (.A1(_07227_),
    .A2(_07245_),
    .Z(_07246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15286_ (.A1(\filters.high[12] ),
    .A2(_07085_),
    .B(_07086_),
    .ZN(_07247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15287_ (.A1(_07058_),
    .A2(_07246_),
    .B(_07247_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15288_ (.A1(_05779_),
    .A2(_07243_),
    .B(_07241_),
    .ZN(_07248_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15289_ (.A1(_01782_),
    .A2(_02068_),
    .A3(_07238_),
    .ZN(_07249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15290_ (.A1(_07236_),
    .A2(_07237_),
    .B(_07249_),
    .ZN(_07250_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15291_ (.A1(_07234_),
    .A2(_07239_),
    .Z(_07251_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15292_ (.A1(_07234_),
    .A2(_07239_),
    .Z(_07252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15293_ (.A1(_07230_),
    .A2(_07251_),
    .B(_07252_),
    .ZN(_07253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15294_ (.A1(_07250_),
    .A2(_07253_),
    .Z(_07254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15295_ (.A1(\filters.low[13] ),
    .A2(_07254_),
    .Z(_07255_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15296_ (.I(_07255_),
    .ZN(_07256_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _15297_ (.A1(_05876_),
    .A2(_05878_),
    .A3(_07256_),
    .Z(_07257_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15298_ (.A1(_07248_),
    .A2(_07257_),
    .ZN(_07258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15299_ (.A1(_05780_),
    .A2(_07243_),
    .ZN(_07259_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15300_ (.A1(_05779_),
    .A2(_07243_),
    .Z(_07260_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _15301_ (.A1(_07259_),
    .A2(_07260_),
    .A3(_07244_),
    .Z(_07261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15302_ (.A1(_07226_),
    .A2(_07245_),
    .B(_07261_),
    .ZN(_07262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15303_ (.A1(_07258_),
    .A2(_07262_),
    .B(_07052_),
    .ZN(_07263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15304_ (.A1(_07258_),
    .A2(_07262_),
    .B(_07263_),
    .ZN(_07264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15305_ (.A1(\filters.high[13] ),
    .A2(_07055_),
    .B(_06914_),
    .ZN(_07265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15306_ (.A1(_07264_),
    .A2(_07265_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15307_ (.A1(_07250_),
    .A2(_07253_),
    .Z(_07266_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15308_ (.A1(\filters.low[14] ),
    .A2(_07266_),
    .Z(_07267_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15309_ (.A1(_05993_),
    .A2(_07267_),
    .Z(_07268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15310_ (.A1(_03441_),
    .A2(_07254_),
    .ZN(_07269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15311_ (.I(_07269_),
    .ZN(_07270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15312_ (.A1(_05879_),
    .A2(_07256_),
    .B(_07270_),
    .ZN(_07271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15313_ (.A1(_07268_),
    .A2(_07271_),
    .Z(_07272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15314_ (.A1(_07245_),
    .A2(_07258_),
    .ZN(_07273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15315_ (.A1(_07241_),
    .A2(_07260_),
    .B(_07257_),
    .ZN(_07274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15316_ (.A1(_07241_),
    .A2(_07260_),
    .A3(_07257_),
    .ZN(_07275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15317_ (.A1(_07261_),
    .A2(_07274_),
    .B(_07275_),
    .ZN(_07276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15318_ (.A1(_07227_),
    .A2(_07273_),
    .B(_07276_),
    .ZN(_07277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15319_ (.A1(_07272_),
    .A2(_07277_),
    .Z(_07278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15320_ (.A1(_07272_),
    .A2(_07277_),
    .B(_07004_),
    .ZN(_07279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15321_ (.A1(_07278_),
    .A2(_07279_),
    .ZN(_07280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15322_ (.A1(\filters.high[14] ),
    .A2(_06979_),
    .B(_07280_),
    .ZN(_07281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15323_ (.A1(_06942_),
    .A2(_07281_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _15324_ (.A1(\filters.low[15] ),
    .A2(_06090_),
    .ZN(_07282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15325_ (.A1(_05993_),
    .A2(_07267_),
    .ZN(_07283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15326_ (.A1(_03457_),
    .A2(_07266_),
    .B(_07283_),
    .ZN(_07284_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15327_ (.A1(_07282_),
    .A2(_07284_),
    .Z(_07285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _15328_ (.A1(_07282_),
    .A2(_07284_),
    .ZN(_07286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15329_ (.A1(_07285_),
    .A2(_07286_),
    .ZN(_07287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15330_ (.A1(_07268_),
    .A2(_07271_),
    .B(_07278_),
    .ZN(_07288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15331_ (.A1(_07287_),
    .A2(_07288_),
    .B(_07110_),
    .ZN(_07289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15332_ (.A1(_07287_),
    .A2(_07288_),
    .B(_07289_),
    .ZN(_07290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15333_ (.A1(_03469_),
    .A2(_06934_),
    .B(_07290_),
    .C(_07219_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15334_ (.A1(_07221_),
    .A2(_07225_),
    .B(_07273_),
    .ZN(_07291_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _15335_ (.A1(_07268_),
    .A2(_07271_),
    .ZN(_07292_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _15336_ (.A1(_07292_),
    .A2(_07285_),
    .A3(_07286_),
    .ZN(_07293_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _15337_ (.A1(_07292_),
    .A2(_07276_),
    .A3(_07285_),
    .A4(_07286_),
    .ZN(_07294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15338_ (.A1(_07268_),
    .A2(_07271_),
    .ZN(_07295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15339_ (.A1(_07282_),
    .A2(_07284_),
    .ZN(_07296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15340_ (.A1(_07295_),
    .A2(_07286_),
    .B(_07296_),
    .ZN(_07297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _15341_ (.A1(_07291_),
    .A2(_07293_),
    .B(_07294_),
    .C(_07297_),
    .ZN(_07298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15342_ (.A1(_03470_),
    .A2(_06090_),
    .ZN(_07299_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15343_ (.A1(\filters.low[16] ),
    .A2(_06201_),
    .ZN(_07300_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15344_ (.A1(_07299_),
    .A2(_07300_),
    .ZN(_07301_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15345_ (.A1(_07298_),
    .A2(_07301_),
    .ZN(_07302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15346_ (.A1(\filters.high[16] ),
    .A2(_07085_),
    .B(_07086_),
    .ZN(_07303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15347_ (.A1(_07058_),
    .A2(_07302_),
    .B(_07303_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15348_ (.A1(\filters.low[16] ),
    .A2(_06311_),
    .Z(_07304_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _15349_ (.A1(\filters.low[17] ),
    .A2(_06317_),
    .A3(_07304_),
    .ZN(_07305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15350_ (.A1(_07299_),
    .A2(_07300_),
    .ZN(_07306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15351_ (.A1(_07298_),
    .A2(_07301_),
    .B(_07306_),
    .ZN(_07307_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15352_ (.A1(_07305_),
    .A2(_07307_),
    .ZN(_07308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15353_ (.A1(_06943_),
    .A2(_07308_),
    .ZN(_07309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15354_ (.I(_06826_),
    .Z(_07310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15355_ (.A1(\filters.high[17] ),
    .A2(_07055_),
    .B(_07310_),
    .ZN(_07311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15356_ (.A1(_07309_),
    .A2(_07311_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15357_ (.A1(\filters.high[18] ),
    .A2(_06979_),
    .ZN(_07312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15358_ (.A1(\filters.low[17] ),
    .A2(_06317_),
    .ZN(_07313_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15359_ (.A1(\filters.low[18] ),
    .A2(_06419_),
    .Z(_07314_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15360_ (.A1(_07313_),
    .A2(_07314_),
    .Z(_07315_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15361_ (.A1(_07301_),
    .A2(_07305_),
    .Z(_07316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15362_ (.I(\filters.low[17] ),
    .Z(_07317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15363_ (.A1(_07317_),
    .A2(_06318_),
    .Z(_07318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15364_ (.A1(_07304_),
    .A2(_07318_),
    .ZN(_07319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15365_ (.A1(_07304_),
    .A2(_07318_),
    .B(_07306_),
    .ZN(_07320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15366_ (.A1(_07319_),
    .A2(_07320_),
    .ZN(_07321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15367_ (.A1(_07298_),
    .A2(_07316_),
    .B(_07321_),
    .ZN(_07322_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15368_ (.A1(_07315_),
    .A2(_07322_),
    .ZN(_07323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15369_ (.A1(_07005_),
    .A2(_07323_),
    .ZN(_07324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15370_ (.A1(_07312_),
    .A2(_07324_),
    .B(_03750_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15371_ (.A1(\filters.low[18] ),
    .A2(_06419_),
    .Z(_07325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15372_ (.A1(\filters.low[19] ),
    .A2(_06521_),
    .Z(_07326_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15373_ (.A1(_07325_),
    .A2(_07326_),
    .ZN(_07327_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15374_ (.A1(_07317_),
    .A2(_06318_),
    .A3(_07314_),
    .ZN(_07328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15375_ (.A1(_07317_),
    .A2(_06318_),
    .B(_07314_),
    .ZN(_07329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15376_ (.A1(_07328_),
    .A2(_07322_),
    .B(_07329_),
    .ZN(_07330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15377_ (.A1(_07327_),
    .A2(_07330_),
    .ZN(_07331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15378_ (.I(_07004_),
    .Z(_07332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15379_ (.A1(\filters.high[19] ),
    .A2(_07332_),
    .B(_07086_),
    .ZN(_07333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15380_ (.A1(_07058_),
    .A2(_07331_),
    .B(_07333_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15381_ (.I(_07057_),
    .Z(_07334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15382_ (.A1(\filters.low[19] ),
    .A2(_06522_),
    .ZN(_07335_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15383_ (.A1(\filters.low[20] ),
    .A2(_06625_),
    .ZN(_07336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15384_ (.A1(_07335_),
    .A2(_07336_),
    .Z(_07337_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15385_ (.A1(_07315_),
    .A2(_07327_),
    .Z(_07338_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _15386_ (.A1(_07315_),
    .A2(_07316_),
    .A3(_07327_),
    .Z(_07339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15387_ (.A1(_07325_),
    .A2(_07326_),
    .ZN(_07340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15388_ (.A1(_07325_),
    .A2(_07326_),
    .ZN(_07341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15389_ (.A1(_07329_),
    .A2(_07340_),
    .B(_07341_),
    .ZN(_07342_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _15390_ (.A1(_07321_),
    .A2(_07338_),
    .B1(_07339_),
    .B2(_07298_),
    .C(_07342_),
    .ZN(_07343_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15391_ (.A1(_07337_),
    .A2(_07343_),
    .ZN(_07344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15392_ (.I(_06738_),
    .Z(_07345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15393_ (.A1(\filters.high[20] ),
    .A2(_07332_),
    .B(_07345_),
    .ZN(_07346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15394_ (.A1(_07334_),
    .A2(_07344_),
    .B(_07346_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15395_ (.A1(_07335_),
    .A2(_07336_),
    .ZN(_07347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15396_ (.A1(_07337_),
    .A2(_07343_),
    .ZN(_07348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15397_ (.A1(_07347_),
    .A2(_07348_),
    .ZN(_07349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15398_ (.I(\filters.low[21] ),
    .Z(_07350_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15399_ (.A1(\filters.low[20] ),
    .A2(_06625_),
    .Z(_07351_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _15400_ (.A1(_07350_),
    .A2(_06780_),
    .A3(_07351_),
    .Z(_07352_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15401_ (.A1(_07349_),
    .A2(_07352_),
    .ZN(_07353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15402_ (.A1(\filters.high[21] ),
    .A2(_07332_),
    .B(_07345_),
    .ZN(_07354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15403_ (.A1(_07334_),
    .A2(_07353_),
    .B(_07354_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15404_ (.A1(\filters.high[22] ),
    .A2(_06943_),
    .ZN(_07355_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15405_ (.A1(_07350_),
    .A2(_06741_),
    .Z(_07356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15406_ (.A1(\filters.low[22] ),
    .A2(_06800_),
    .Z(_07357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _15407_ (.A1(_07356_),
    .A2(_07357_),
    .Z(_07358_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _15408_ (.A1(_07337_),
    .A2(_07352_),
    .Z(_07359_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15409_ (.A1(_07350_),
    .A2(_06860_),
    .Z(_07360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15410_ (.A1(_07351_),
    .A2(_07360_),
    .ZN(_07361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15411_ (.A1(_07351_),
    .A2(_07360_),
    .B(_07347_),
    .ZN(_07362_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15412_ (.A1(_07361_),
    .A2(_07362_),
    .Z(_07363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15413_ (.A1(_07343_),
    .A2(_07359_),
    .B(_07363_),
    .ZN(_07364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15414_ (.I(_07364_),
    .ZN(_07365_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15415_ (.A1(_07358_),
    .A2(_07365_),
    .Z(_07366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15416_ (.A1(_07085_),
    .A2(_07366_),
    .ZN(_07367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15417_ (.I(_03651_),
    .Z(_07368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15418_ (.A1(_07355_),
    .A2(_07367_),
    .B(_07368_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15419_ (.A1(_07356_),
    .A2(_07357_),
    .ZN(_07369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15420_ (.A1(_07358_),
    .A2(_07365_),
    .B(_07369_),
    .ZN(_07370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15421_ (.A1(\filters.low[22] ),
    .A2(_06860_),
    .ZN(_07371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15422_ (.A1(\filters.low[23] ),
    .A2(_06780_),
    .Z(_07372_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15423_ (.A1(_07371_),
    .A2(_07372_),
    .ZN(_07373_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15424_ (.A1(_07370_),
    .A2(_07373_),
    .Z(_07374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15425_ (.A1(\filters.high[23] ),
    .A2(_07332_),
    .B(_07345_),
    .ZN(_07375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15426_ (.A1(_07334_),
    .A2(_07374_),
    .B(_07375_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15427_ (.A1(_07358_),
    .A2(_07373_),
    .Z(_07376_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _15428_ (.A1(_07358_),
    .A2(_07359_),
    .A3(_07373_),
    .Z(_07377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15429_ (.I(_07371_),
    .ZN(_07378_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _15430_ (.A1(_06846_),
    .A2(_07356_),
    .A3(_07357_),
    .B1(_07372_),
    .B2(_07378_),
    .ZN(_07379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _15431_ (.A1(_07363_),
    .A2(_07376_),
    .B1(_07377_),
    .B2(_07343_),
    .C(_07379_),
    .ZN(_07380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15432_ (.I(\filters.low[24] ),
    .Z(_07381_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15433_ (.A1(_07381_),
    .A2(_06877_),
    .Z(_07382_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _15434_ (.A1(\filters.low[23] ),
    .A2(_06886_),
    .Z(_07383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _15435_ (.I0(_07382_),
    .I1(_07381_),
    .S(_07383_),
    .Z(_07384_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15436_ (.A1(net29),
    .A2(_07384_),
    .Z(_07385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15437_ (.A1(\filters.high[24] ),
    .A2(_07057_),
    .B(_07345_),
    .ZN(_07386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15438_ (.A1(_07334_),
    .A2(_07385_),
    .B(_07386_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15439_ (.I(\filters.high[25] ),
    .ZN(_07387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _15440_ (.A1(_07383_),
    .A2(_07382_),
    .ZN(_07388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _15441_ (.A1(_06861_),
    .A2(_07383_),
    .B(_07380_),
    .C(_07388_),
    .ZN(_07389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15442_ (.I(\filters.low[25] ),
    .Z(_07390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15443_ (.I(_07390_),
    .Z(_07391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15444_ (.A1(_07381_),
    .A2(_06886_),
    .ZN(_07392_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15445_ (.A1(_07390_),
    .A2(_06877_),
    .Z(_07393_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15446_ (.I(_07393_),
    .ZN(_07394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15447_ (.A1(_07392_),
    .A2(_07394_),
    .ZN(_07395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15448_ (.A1(_07391_),
    .A2(_07392_),
    .B(_07395_),
    .ZN(_07396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15449_ (.A1(_07388_),
    .A2(_07389_),
    .B(_07396_),
    .ZN(_07397_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _15450_ (.A1(_07388_),
    .A2(_07389_),
    .A3(_07396_),
    .ZN(_07398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15451_ (.A1(_06958_),
    .A2(_07398_),
    .ZN(_07399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _15452_ (.A1(_07387_),
    .A2(_06934_),
    .B1(_07397_),
    .B2(_07399_),
    .C(_06941_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15453_ (.I(_01944_),
    .Z(_07400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15454_ (.I(\filters.low[26] ),
    .Z(_07401_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15455_ (.A1(\filters.low[26] ),
    .A2(_06877_),
    .Z(_07402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15456_ (.A1(_07390_),
    .A2(_06789_),
    .ZN(_07403_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _15457_ (.I0(_07401_),
    .I1(_07402_),
    .S(_07403_),
    .Z(_07404_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _15458_ (.I0(_07390_),
    .I1(_07393_),
    .S(_07392_),
    .Z(_07405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15459_ (.A1(_07384_),
    .A2(_07405_),
    .ZN(_07406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _15460_ (.A1(_07391_),
    .A2(_07388_),
    .B1(_07394_),
    .B2(_07392_),
    .ZN(_07407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15461_ (.A1(net50),
    .A2(_07406_),
    .B(_07407_),
    .ZN(_07408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15462_ (.A1(_07404_),
    .A2(_07408_),
    .ZN(_07409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15463_ (.A1(_07404_),
    .A2(_07408_),
    .ZN(_07410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15464_ (.A1(_06933_),
    .A2(_07410_),
    .ZN(_07411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15465_ (.A1(\filters.high[26] ),
    .A2(_06958_),
    .B1(_07409_),
    .B2(_07411_),
    .ZN(_07412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15466_ (.A1(_07400_),
    .A2(_07412_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15467_ (.I(\filters.low[27] ),
    .Z(_07413_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15468_ (.A1(\filters.low[27] ),
    .A2(_06886_),
    .Z(_07414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15469_ (.A1(_07401_),
    .A2(_06759_),
    .ZN(_07415_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _15470_ (.I0(_07413_),
    .I1(_07414_),
    .S(_07415_),
    .Z(_07416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15471_ (.A1(_07391_),
    .A2(_06791_),
    .B(_07402_),
    .ZN(_07417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15472_ (.A1(_07404_),
    .A2(_07408_),
    .B(_07417_),
    .ZN(_07418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15473_ (.A1(_07416_),
    .A2(_07418_),
    .B(_07052_),
    .ZN(_07419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15474_ (.A1(_07416_),
    .A2(_07418_),
    .B(_07419_),
    .ZN(_07420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15475_ (.A1(\filters.high[27] ),
    .A2(_07005_),
    .B(_07310_),
    .ZN(_07421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15476_ (.A1(_07420_),
    .A2(_07421_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15477_ (.A1(_07404_),
    .A2(_07416_),
    .ZN(_07422_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15478_ (.A1(_07406_),
    .A2(_07422_),
    .Z(_07423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15479_ (.A1(_07401_),
    .A2(_06791_),
    .B(_07414_),
    .ZN(_07424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15480_ (.A1(_07413_),
    .A2(_07417_),
    .B(_07424_),
    .ZN(_07425_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _15481_ (.A1(_07407_),
    .A2(_07422_),
    .B1(_07423_),
    .B2(_07380_),
    .C(_07425_),
    .ZN(_07426_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15482_ (.A1(_07413_),
    .A2(_06790_),
    .Z(_07427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15483_ (.A1(\filters.low[28] ),
    .A2(_06742_),
    .Z(_07428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15484_ (.A1(_07427_),
    .A2(_07428_),
    .ZN(_07429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15485_ (.A1(_06899_),
    .A2(_07427_),
    .B(_07429_),
    .ZN(_07430_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15486_ (.A1(_07426_),
    .A2(_07430_),
    .ZN(_07431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15487_ (.I(_06738_),
    .Z(_07432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15488_ (.A1(\filters.high[28] ),
    .A2(_07057_),
    .B(_07432_),
    .ZN(_07433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15489_ (.A1(_07055_),
    .A2(_07431_),
    .B(_07433_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15490_ (.A1(\filters.low[28] ),
    .A2(_06790_),
    .Z(_07434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15491_ (.I(\filters.low[29] ),
    .Z(_07435_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15492_ (.A1(_07435_),
    .A2(_06742_),
    .Z(_07436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15493_ (.A1(_07434_),
    .A2(_07436_),
    .ZN(_07437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15494_ (.A1(_06906_),
    .A2(_07434_),
    .B(_07437_),
    .ZN(_07438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15495_ (.A1(_07426_),
    .A2(_07430_),
    .B(_07429_),
    .ZN(_07439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15496_ (.A1(_07438_),
    .A2(_07439_),
    .B(_07052_),
    .ZN(_07440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15497_ (.A1(_07438_),
    .A2(_07439_),
    .B(_07440_),
    .ZN(_07441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15498_ (.A1(\filters.high[29] ),
    .A2(_07005_),
    .B(_07310_),
    .ZN(_07442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15499_ (.A1(_07441_),
    .A2(_07442_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15500_ (.A1(\filters.high[30] ),
    .A2(_06943_),
    .ZN(_07443_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15501_ (.A1(_07430_),
    .A2(_07438_),
    .Z(_07444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _15502_ (.A1(_07435_),
    .A2(_07429_),
    .B1(_07444_),
    .B2(_07426_),
    .C(_07437_),
    .ZN(_07445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15503_ (.A1(_06916_),
    .A2(_06791_),
    .ZN(_07446_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15504_ (.I(_07446_),
    .ZN(_07447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15505_ (.A1(_06916_),
    .A2(_06744_),
    .ZN(_07448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _15506_ (.A1(_07435_),
    .A2(_06792_),
    .B(_07448_),
    .C(_07447_),
    .ZN(_07449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15507_ (.A1(_07435_),
    .A2(_07447_),
    .B(_07449_),
    .ZN(_07450_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15508_ (.I(_07450_),
    .ZN(_07451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15509_ (.A1(_07445_),
    .A2(_07451_),
    .B(_06976_),
    .ZN(_07452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15510_ (.A1(_07445_),
    .A2(_07451_),
    .B(_07452_),
    .ZN(_07453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15511_ (.A1(_07443_),
    .A2(_07453_),
    .B(_07368_),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15512_ (.I(\filters.high[31] ),
    .ZN(_07454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15513_ (.A1(_07445_),
    .A2(_07451_),
    .ZN(_07455_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _15514_ (.A1(_07449_),
    .A2(_07455_),
    .Z(_07456_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15515_ (.A1(\filters.low[31] ),
    .A2(_07447_),
    .Z(_07457_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15516_ (.I(_07457_),
    .ZN(_07458_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15517_ (.A1(_07456_),
    .A2(_07458_),
    .Z(_07459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15518_ (.A1(_07456_),
    .A2(_07458_),
    .B(_06937_),
    .ZN(_07460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _15519_ (.A1(_07454_),
    .A2(_06934_),
    .B1(_07459_),
    .B2(_07460_),
    .C(_06941_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15520_ (.I(_03204_),
    .Z(_07461_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15521_ (.A1(\filters.mode_vol[7] ),
    .A2(_01783_),
    .B(_03216_),
    .C(_03217_),
    .ZN(_07462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _15522_ (.A1(_01758_),
    .A2(_03430_),
    .B1(_03478_),
    .B2(_01772_),
    .C1(_07461_),
    .C2(_03239_),
    .ZN(_07463_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _15523_ (.A1(_07461_),
    .A2(_07462_),
    .B(_07463_),
    .C(_03757_),
    .ZN(_07464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15524_ (.I(_07464_),
    .Z(_07465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15525_ (.I(_07465_),
    .Z(_07466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15526_ (.A1(_03196_),
    .A2(_04242_),
    .B(_07464_),
    .ZN(_07467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15527_ (.I(_07467_),
    .Z(_07468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15528_ (.I(_07468_),
    .Z(_07469_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _15529_ (.A1(_03204_),
    .A2(_03206_),
    .A3(_03217_),
    .ZN(_07470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15530_ (.I(_07470_),
    .Z(_07471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15531_ (.A1(\channels.sample3[0] ),
    .A2(_07471_),
    .ZN(_07472_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15532_ (.A1(_03265_),
    .A2(_07471_),
    .B(_07472_),
    .C(_03221_),
    .ZN(_07473_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15533_ (.A1(\channels.sample2[0] ),
    .A2(_06091_),
    .B(_07473_),
    .C(_03346_),
    .ZN(_07474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15534_ (.A1(\channels.sample1[0] ),
    .A2(_03402_),
    .ZN(_07475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15535_ (.A1(_07474_),
    .A2(_07475_),
    .ZN(_07476_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15536_ (.A1(\filters.sample_buff[0] ),
    .A2(_07476_),
    .Z(_07477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15537_ (.A1(\filters.sample_buff[0] ),
    .A2(_07466_),
    .B1(_07469_),
    .B2(_07477_),
    .ZN(_07478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15538_ (.A1(_07400_),
    .A2(_07478_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15539_ (.I(_07464_),
    .Z(_07479_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15540_ (.A1(\filters.sample_buff[0] ),
    .A2(_07476_),
    .Z(_07480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15541_ (.I(_07470_),
    .Z(_07481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15542_ (.A1(\channels.sample3[1] ),
    .A2(_07470_),
    .ZN(_07482_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15543_ (.A1(_03266_),
    .A2(_07481_),
    .B(_07482_),
    .C(_03220_),
    .ZN(_07483_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15544_ (.A1(\channels.sample2[1] ),
    .A2(_03221_),
    .B(_07483_),
    .C(_03231_),
    .ZN(_07484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15545_ (.A1(\channels.sample1[1] ),
    .A2(_03337_),
    .ZN(_07485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15546_ (.A1(_07484_),
    .A2(_07485_),
    .ZN(_07486_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15547_ (.A1(\filters.sample_buff[1] ),
    .A2(_07486_),
    .Z(_07487_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15548_ (.A1(_07480_),
    .A2(_07487_),
    .Z(_07488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15549_ (.A1(\filters.sample_buff[1] ),
    .A2(_07479_),
    .B1(_07469_),
    .B2(_07488_),
    .ZN(_07489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15550_ (.A1(_07400_),
    .A2(_07489_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15551_ (.A1(\filters.sample_buff[1] ),
    .A2(_07486_),
    .ZN(_07490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15552_ (.A1(_07480_),
    .A2(_07487_),
    .ZN(_07491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15553_ (.A1(\channels.sample3[2] ),
    .A2(_07481_),
    .ZN(_07492_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15554_ (.A1(_03283_),
    .A2(_07481_),
    .B(_07492_),
    .C(_03377_),
    .ZN(_07493_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15555_ (.A1(\channels.sample2[2] ),
    .A2(_03348_),
    .B(_07493_),
    .C(_03231_),
    .ZN(_07494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15556_ (.A1(\channels.sample1[2] ),
    .A2(_03337_),
    .ZN(_07495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15557_ (.A1(_07494_),
    .A2(_07495_),
    .ZN(_07496_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15558_ (.A1(\filters.sample_buff[2] ),
    .A2(_07496_),
    .ZN(_07497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15559_ (.A1(_07490_),
    .A2(_07491_),
    .B(_07497_),
    .ZN(_07498_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15560_ (.A1(_07490_),
    .A2(_07491_),
    .A3(_07497_),
    .Z(_07499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15561_ (.A1(_07498_),
    .A2(_07499_),
    .ZN(_07500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15562_ (.A1(\filters.sample_buff[2] ),
    .A2(_07479_),
    .B1(_07469_),
    .B2(_07500_),
    .ZN(_07501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15563_ (.A1(_07400_),
    .A2(_07501_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15564_ (.I(_07464_),
    .Z(_07502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15565_ (.A1(\filters.sample_buff[3] ),
    .A2(_07502_),
    .ZN(_07503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15566_ (.I(_07467_),
    .Z(_07504_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15567_ (.A1(\filters.sample_buff[2] ),
    .A2(_07496_),
    .Z(_07505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15568_ (.I(_07481_),
    .Z(_07506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15569_ (.A1(\channels.sample3[3] ),
    .A2(_07471_),
    .ZN(_07507_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15570_ (.A1(_03299_),
    .A2(_07506_),
    .B(_07507_),
    .C(_03378_),
    .ZN(_07508_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15571_ (.A1(\channels.sample2[3] ),
    .A2(_03222_),
    .B(_07508_),
    .C(_03346_),
    .ZN(_07509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15572_ (.A1(\channels.sample1[3] ),
    .A2(_03402_),
    .ZN(_07510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15573_ (.A1(_07509_),
    .A2(_07510_),
    .ZN(_07511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15574_ (.A1(\filters.sample_buff[3] ),
    .A2(_07511_),
    .Z(_07512_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15575_ (.A1(_07505_),
    .A2(_07498_),
    .A3(_07512_),
    .Z(_07513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15576_ (.A1(_07505_),
    .A2(_07498_),
    .B(_07512_),
    .ZN(_07514_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15577_ (.A1(_07504_),
    .A2(_07513_),
    .A3(_07514_),
    .ZN(_07515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15578_ (.A1(_07503_),
    .A2(_07515_),
    .B(_07368_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15579_ (.I(_01944_),
    .Z(_07516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15580_ (.A1(\filters.sample_buff[3] ),
    .A2(_07511_),
    .ZN(_07517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15581_ (.A1(\channels.sample3[4] ),
    .A2(_07471_),
    .ZN(_07518_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15582_ (.A1(_03311_),
    .A2(_07506_),
    .B(_07518_),
    .C(_06091_),
    .ZN(_07519_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15583_ (.A1(\channels.sample2[4] ),
    .A2(_03379_),
    .B(_07519_),
    .C(_03232_),
    .ZN(_07520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15584_ (.A1(\channels.sample1[4] ),
    .A2(_03402_),
    .ZN(_07521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15585_ (.A1(_07520_),
    .A2(_07521_),
    .ZN(_07522_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15586_ (.A1(\filters.sample_buff[4] ),
    .A2(_07522_),
    .Z(_07523_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15587_ (.I(_07523_),
    .ZN(_07524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15588_ (.A1(_07517_),
    .A2(_07514_),
    .B(_07524_),
    .ZN(_07525_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15589_ (.A1(_07517_),
    .A2(_07514_),
    .A3(_07524_),
    .Z(_07526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15590_ (.A1(_07525_),
    .A2(_07526_),
    .ZN(_07527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15591_ (.A1(\filters.sample_buff[4] ),
    .A2(_07479_),
    .B1(_07469_),
    .B2(_07527_),
    .ZN(_07528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15592_ (.A1(_07516_),
    .A2(_07528_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15593_ (.A1(\filters.sample_buff[5] ),
    .A2(_07502_),
    .ZN(_07529_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15594_ (.A1(\filters.sample_buff[4] ),
    .A2(_07522_),
    .Z(_07530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15595_ (.I(_07506_),
    .Z(_07531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15596_ (.A1(_01939_),
    .A2(_07506_),
    .ZN(_07532_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15597_ (.A1(_03328_),
    .A2(_07531_),
    .B(_07532_),
    .C(_06092_),
    .ZN(_07533_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15598_ (.A1(\channels.sample2[5] ),
    .A2(_03380_),
    .B(_07533_),
    .C(_03233_),
    .ZN(_07534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15599_ (.A1(\channels.sample1[5] ),
    .A2(_03403_),
    .ZN(_07535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15600_ (.A1(_07534_),
    .A2(_07535_),
    .ZN(_07536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15601_ (.A1(\filters.sample_buff[5] ),
    .A2(_07536_),
    .Z(_07537_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15602_ (.A1(_07530_),
    .A2(_07525_),
    .A3(_07537_),
    .Z(_07538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15603_ (.A1(_07530_),
    .A2(_07525_),
    .B(_07537_),
    .ZN(_07539_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15604_ (.A1(_07504_),
    .A2(_07538_),
    .A3(_07539_),
    .ZN(_07540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15605_ (.A1(_07529_),
    .A2(_07540_),
    .B(_07368_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15606_ (.I(_07467_),
    .Z(_07541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15607_ (.A1(\filters.sample_buff[5] ),
    .A2(_07536_),
    .ZN(_07542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15608_ (.A1(\channels.sample3[6] ),
    .A2(_07531_),
    .ZN(_07543_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15609_ (.A1(_03344_),
    .A2(_07531_),
    .B(_07543_),
    .C(_06202_),
    .ZN(_07544_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15610_ (.A1(\channels.sample2[6] ),
    .A2(_06420_),
    .B(_07544_),
    .C(_03233_),
    .ZN(_07545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15611_ (.A1(\channels.sample1[6] ),
    .A2(_03403_),
    .ZN(_07546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15612_ (.A1(_07545_),
    .A2(_07546_),
    .ZN(_07547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15613_ (.A1(\filters.sample_buff[6] ),
    .A2(_07547_),
    .Z(_07548_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15614_ (.I(_07548_),
    .ZN(_07549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15615_ (.A1(_07542_),
    .A2(_07539_),
    .B(_07549_),
    .ZN(_07550_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15616_ (.A1(_07542_),
    .A2(_07539_),
    .A3(_07549_),
    .Z(_07551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15617_ (.A1(_07550_),
    .A2(_07551_),
    .ZN(_07552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15618_ (.A1(\filters.sample_buff[6] ),
    .A2(_07479_),
    .B1(_07541_),
    .B2(_07552_),
    .ZN(_07553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15619_ (.A1(_07516_),
    .A2(_07553_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15620_ (.A1(\filters.sample_buff[7] ),
    .A2(_07502_),
    .ZN(_07554_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15621_ (.A1(\filters.sample_buff[6] ),
    .A2(_07547_),
    .Z(_07555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15622_ (.I(_07531_),
    .Z(_07556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15623_ (.A1(_01989_),
    .A2(_07556_),
    .ZN(_07557_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15624_ (.A1(_03360_),
    .A2(_07556_),
    .B(_07557_),
    .C(_06733_),
    .ZN(_07558_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15625_ (.A1(\channels.sample2[7] ),
    .A2(_03397_),
    .B(_07558_),
    .C(_03234_),
    .ZN(_07559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15626_ (.A1(\channels.sample1[7] ),
    .A2(_03429_),
    .ZN(_07560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15627_ (.A1(_07559_),
    .A2(_07560_),
    .ZN(_07561_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15628_ (.A1(\filters.sample_buff[7] ),
    .A2(_07561_),
    .Z(_07562_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15629_ (.A1(_07555_),
    .A2(_07550_),
    .A3(_07562_),
    .Z(_07563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15630_ (.A1(_07555_),
    .A2(_07550_),
    .B(_07562_),
    .ZN(_07564_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15631_ (.A1(_07504_),
    .A2(_07563_),
    .A3(_07564_),
    .ZN(_07565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15632_ (.I(_03650_),
    .Z(_07566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15633_ (.I(_07566_),
    .Z(_07567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15634_ (.A1(_07554_),
    .A2(_07565_),
    .B(_07567_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15635_ (.A1(\filters.sample_buff[7] ),
    .A2(_07561_),
    .ZN(_07568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15636_ (.I(_07556_),
    .Z(_07569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15637_ (.A1(\channels.sample3[8] ),
    .A2(_07556_),
    .ZN(_07570_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15638_ (.A1(_03374_),
    .A2(_07569_),
    .B(_07570_),
    .C(_03397_),
    .ZN(_07571_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _15639_ (.A1(\channels.sample2[8] ),
    .A2(_03225_),
    .B(_07571_),
    .C(_03234_),
    .ZN(_07572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15640_ (.A1(\channels.sample1[8] ),
    .A2(_03429_),
    .ZN(_07573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15641_ (.A1(_07572_),
    .A2(_07573_),
    .ZN(_07574_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15642_ (.A1(\filters.sample_buff[8] ),
    .A2(_07574_),
    .Z(_07575_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15643_ (.I(_07575_),
    .ZN(_07576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15644_ (.A1(_07568_),
    .A2(_07564_),
    .B(_07576_),
    .ZN(_07577_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15645_ (.A1(_07568_),
    .A2(_07564_),
    .A3(_07576_),
    .Z(_07578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15646_ (.A1(_07577_),
    .A2(_07578_),
    .ZN(_07579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15647_ (.A1(\filters.sample_buff[8] ),
    .A2(_07465_),
    .B1(_07541_),
    .B2(_07579_),
    .ZN(_07580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15648_ (.A1(_07516_),
    .A2(_07580_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15649_ (.A1(\filters.sample_buff[9] ),
    .A2(_07466_),
    .ZN(_07581_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15650_ (.A1(\filters.sample_buff[8] ),
    .A2(_07574_),
    .Z(_07582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15651_ (.I(_07569_),
    .Z(_07583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15652_ (.A1(_02040_),
    .A2(_07569_),
    .ZN(_07584_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15653_ (.A1(_03393_),
    .A2(_07583_),
    .B(_07584_),
    .C(_03225_),
    .ZN(_07585_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15654_ (.A1(\channels.sample2[9] ),
    .A2(_03426_),
    .B(_07585_),
    .C(_03235_),
    .ZN(_07586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15655_ (.A1(\channels.sample1[9] ),
    .A2(_03429_),
    .ZN(_07587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15656_ (.A1(_07586_),
    .A2(_07587_),
    .ZN(_07588_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15657_ (.A1(\filters.sample_buff[9] ),
    .A2(_07588_),
    .Z(_07589_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15658_ (.A1(_07582_),
    .A2(_07577_),
    .A3(_07589_),
    .Z(_07590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15659_ (.A1(_07582_),
    .A2(_07577_),
    .B(_07589_),
    .ZN(_07591_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15660_ (.A1(_07504_),
    .A2(_07590_),
    .A3(_07591_),
    .ZN(_07592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15661_ (.A1(_07581_),
    .A2(_07592_),
    .B(_07567_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15662_ (.A1(\filters.sample_buff[9] ),
    .A2(_07588_),
    .ZN(_07593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15663_ (.A1(\channels.sample3[10] ),
    .A2(_07569_),
    .ZN(_07594_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15664_ (.A1(_03411_),
    .A2(_07583_),
    .B(_07594_),
    .C(_03426_),
    .ZN(_07595_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15665_ (.A1(\channels.sample2[10] ),
    .A2(_03426_),
    .B(_07595_),
    .C(_03236_),
    .ZN(_07596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15666_ (.A1(\channels.sample1[10] ),
    .A2(_03430_),
    .ZN(_07597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15667_ (.A1(_07596_),
    .A2(_07597_),
    .ZN(_07598_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15668_ (.A1(\filters.sample_buff[10] ),
    .A2(_07598_),
    .Z(_07599_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15669_ (.I(_07599_),
    .ZN(_07600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15670_ (.A1(_07593_),
    .A2(_07591_),
    .B(_07600_),
    .ZN(_07601_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15671_ (.A1(_07593_),
    .A2(_07591_),
    .A3(_07600_),
    .Z(_07602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15672_ (.A1(_07601_),
    .A2(_07602_),
    .ZN(_07603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15673_ (.A1(\filters.sample_buff[10] ),
    .A2(_07465_),
    .B1(_07541_),
    .B2(_07603_),
    .ZN(_07604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15674_ (.A1(_07516_),
    .A2(_07604_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15675_ (.A1(\filters.sample_buff[11] ),
    .A2(_07466_),
    .ZN(_07605_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15676_ (.A1(\filters.sample_buff[10] ),
    .A2(_07598_),
    .Z(_07606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15677_ (.A1(_02068_),
    .A2(_07583_),
    .ZN(_07607_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15678_ (.A1(_03423_),
    .A2(_07583_),
    .B(_07607_),
    .C(_03226_),
    .ZN(_07608_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15679_ (.A1(\channels.sample2[11] ),
    .A2(_03227_),
    .B(_07608_),
    .C(_03236_),
    .ZN(_07609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15680_ (.A1(\channels.sample1[11] ),
    .A2(_03430_),
    .ZN(_07610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15681_ (.A1(_07609_),
    .A2(_07610_),
    .ZN(_07611_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15682_ (.A1(\filters.sample_buff[11] ),
    .A2(_07611_),
    .Z(_07612_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15683_ (.A1(_07606_),
    .A2(_07601_),
    .A3(_07612_),
    .Z(_07613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15684_ (.A1(_07606_),
    .A2(_07601_),
    .B(_07612_),
    .ZN(_07614_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15685_ (.A1(_07468_),
    .A2(_07613_),
    .A3(_07614_),
    .ZN(_07615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15686_ (.A1(_07605_),
    .A2(_07615_),
    .B(_07567_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15687_ (.I(_01943_),
    .Z(_07616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15688_ (.I(_07616_),
    .Z(_07617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15689_ (.A1(\filters.sample_buff[11] ),
    .A2(_07611_),
    .ZN(_07618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15690_ (.A1(_07618_),
    .A2(_07614_),
    .ZN(_07619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15691_ (.A1(_03241_),
    .A2(_03239_),
    .ZN(_07620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15692_ (.I(_07620_),
    .Z(_07621_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15693_ (.A1(\filters.sample_buff[12] ),
    .A2(_03452_),
    .A3(_07621_),
    .Z(_07622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15694_ (.A1(_03452_),
    .A2(_07621_),
    .B(\filters.sample_buff[12] ),
    .ZN(_07623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15695_ (.A1(_07622_),
    .A2(_07623_),
    .ZN(_07624_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15696_ (.A1(_07619_),
    .A2(_07624_),
    .Z(_07625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15697_ (.A1(\filters.sample_buff[12] ),
    .A2(_07465_),
    .B1(_07541_),
    .B2(_07625_),
    .ZN(_07626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15698_ (.A1(_07617_),
    .A2(_07626_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15699_ (.A1(\filters.sample_buff[13] ),
    .A2(_07466_),
    .ZN(_07627_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15700_ (.A1(_07619_),
    .A2(_07624_),
    .Z(_07628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15701_ (.A1(\filters.sample_filtered[14] ),
    .A2(_07620_),
    .ZN(_07629_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15702_ (.A1(\filters.sample_buff[13] ),
    .A2(_07629_),
    .ZN(_07630_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _15703_ (.A1(_07622_),
    .A2(_07628_),
    .A3(_07630_),
    .Z(_07631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15704_ (.A1(_07622_),
    .A2(_07628_),
    .B(_07630_),
    .ZN(_07632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15705_ (.A1(_07468_),
    .A2(_07631_),
    .A3(_07632_),
    .ZN(_07633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15706_ (.A1(_07627_),
    .A2(_07633_),
    .B(_07567_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15707_ (.I(\filters.sample_buff[14] ),
    .ZN(_07634_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15708_ (.A1(\filters.sample_buff[13] ),
    .A2(_03454_),
    .A3(_07621_),
    .ZN(_07635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15709_ (.A1(\filters.sample_filtered[15] ),
    .A2(_07621_),
    .ZN(_07636_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15710_ (.A1(_07634_),
    .A2(_07636_),
    .Z(_07637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15711_ (.A1(_07635_),
    .A2(_07632_),
    .B(_07637_),
    .ZN(_07638_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15712_ (.A1(_07635_),
    .A2(_07632_),
    .A3(_07637_),
    .ZN(_07639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15713_ (.A1(_07468_),
    .A2(_07639_),
    .ZN(_07640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15714_ (.A1(_07638_),
    .A2(_07640_),
    .ZN(_07641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15715_ (.A1(_07634_),
    .A2(_07502_),
    .B(_07641_),
    .C(_07219_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15716_ (.I(\channels.exp_periods[3][0] ),
    .Z(_07642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15717_ (.I(_07642_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15718_ (.I(\channels.exp_periods[3][1] ),
    .Z(_07643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15719_ (.I(_07643_),
    .Z(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15720_ (.I(\channels.exp_periods[3][2] ),
    .Z(_07644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15721_ (.I(_07644_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15722_ (.I(\channels.exp_periods[3][3] ),
    .Z(_07645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15723_ (.I(_07645_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15724_ (.I(\channels.exp_periods[3][4] ),
    .Z(_07646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15725_ (.I(_07646_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15726_ (.A1(_03218_),
    .A2(_03757_),
    .ZN(_07647_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _15727_ (.A1(_07461_),
    .A2(_03216_),
    .A3(_07647_),
    .ZN(_07648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15728_ (.I(_07648_),
    .Z(_07649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15729_ (.I(_07649_),
    .Z(_07650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15730_ (.I(_07650_),
    .Z(_07651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15731_ (.I(_07649_),
    .Z(_07652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15732_ (.A1(_05561_),
    .A2(_07652_),
    .B(_07432_),
    .ZN(_07653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15733_ (.A1(_05566_),
    .A2(_07651_),
    .B(_07653_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15734_ (.A1(_03218_),
    .A2(_03758_),
    .A3(_03207_),
    .ZN(_07654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15735_ (.I(_07654_),
    .Z(_07655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15736_ (.I(_07655_),
    .Z(_07656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15737_ (.A1(_05680_),
    .A2(_07656_),
    .ZN(_07657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15738_ (.I(_07648_),
    .Z(_07658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15739_ (.I(_07658_),
    .Z(_07659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15740_ (.A1(_05676_),
    .A2(_07659_),
    .B(_07310_),
    .ZN(_07660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15741_ (.A1(_07657_),
    .A2(_07660_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15742_ (.A1(_05787_),
    .A2(_07656_),
    .ZN(_07661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15743_ (.I(_07658_),
    .Z(_07662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15744_ (.I(_03508_),
    .Z(_07663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15745_ (.I(_07663_),
    .Z(_07664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15746_ (.A1(_03270_),
    .A2(_07662_),
    .B(_07664_),
    .ZN(_07665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15747_ (.A1(_07661_),
    .A2(_07665_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15748_ (.A1(_05889_),
    .A2(_07656_),
    .ZN(_07666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15749_ (.A1(_03284_),
    .A2(_07662_),
    .B(_07664_),
    .ZN(_07667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15750_ (.A1(_07666_),
    .A2(_07667_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15751_ (.A1(_05994_),
    .A2(_07652_),
    .B(_07432_),
    .ZN(_07668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15752_ (.A1(_05998_),
    .A2(_07651_),
    .B(_07668_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15753_ (.A1(_06103_),
    .A2(_07656_),
    .ZN(_07669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15754_ (.A1(_03312_),
    .A2(_07662_),
    .B(_07664_),
    .ZN(_07670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15755_ (.A1(_07669_),
    .A2(_07670_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15756_ (.I(_07655_),
    .Z(_07671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15757_ (.A1(_06209_),
    .A2(_07671_),
    .ZN(_07672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15758_ (.A1(_03331_),
    .A2(_07662_),
    .B(_07664_),
    .ZN(_07673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15759_ (.A1(_07672_),
    .A2(_07673_),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15760_ (.A1(_06315_),
    .A2(_07671_),
    .ZN(_07674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15761_ (.I(_07658_),
    .Z(_07675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15762_ (.I(_07663_),
    .Z(_07676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15763_ (.A1(_03347_),
    .A2(_07675_),
    .B(_07676_),
    .ZN(_07677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15764_ (.A1(_07674_),
    .A2(_07677_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15765_ (.A1(_06424_),
    .A2(_07671_),
    .ZN(_07678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15766_ (.A1(_03362_),
    .A2(_07675_),
    .B(_07676_),
    .ZN(_07679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15767_ (.A1(_07678_),
    .A2(_07679_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15768_ (.A1(_06529_),
    .A2(_07671_),
    .ZN(_07680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15769_ (.A1(_03376_),
    .A2(_07675_),
    .B(_07676_),
    .ZN(_07681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15770_ (.A1(_07680_),
    .A2(_07681_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15771_ (.I(_07654_),
    .Z(_07682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15772_ (.I(_07682_),
    .Z(_07683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15773_ (.A1(_06634_),
    .A2(_07683_),
    .ZN(_07684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15774_ (.A1(_03396_),
    .A2(_07675_),
    .B(_07676_),
    .ZN(_07685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15775_ (.A1(_07684_),
    .A2(_07685_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15776_ (.A1(_03413_),
    .A2(_07652_),
    .B(_07432_),
    .ZN(_07686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15777_ (.A1(_06718_),
    .A2(_07651_),
    .B(_07686_),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15778_ (.I(_03674_),
    .Z(_07687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15779_ (.I(_07687_),
    .Z(_07688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15780_ (.A1(_03424_),
    .A2(_07652_),
    .B(_07688_),
    .ZN(_07689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15781_ (.A1(_06737_),
    .A2(_07651_),
    .B(_07689_),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15782_ (.A1(_06753_),
    .A2(_07683_),
    .ZN(_07690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15783_ (.I(_07658_),
    .Z(_07691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15784_ (.I(_07663_),
    .Z(_07692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15785_ (.A1(_03441_),
    .A2(_07691_),
    .B(_07692_),
    .ZN(_07693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15786_ (.A1(_07690_),
    .A2(_07693_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15787_ (.A1(_06762_),
    .A2(_07683_),
    .ZN(_07694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15788_ (.A1(_03457_),
    .A2(_07691_),
    .B(_07692_),
    .ZN(_07695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15789_ (.A1(_07694_),
    .A2(_07695_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15790_ (.A1(_06771_),
    .A2(_07683_),
    .ZN(_07696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15791_ (.A1(_03470_),
    .A2(_07691_),
    .B(_07692_),
    .ZN(_07697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15792_ (.A1(_07696_),
    .A2(_07697_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15793_ (.I(_07682_),
    .Z(_07698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15794_ (.A1(_06784_),
    .A2(_07698_),
    .ZN(_07699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15795_ (.A1(\filters.low[16] ),
    .A2(_07691_),
    .B(_07692_),
    .ZN(_07700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15796_ (.A1(_07699_),
    .A2(_07700_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15797_ (.A1(_07317_),
    .A2(_07650_),
    .B(_07688_),
    .ZN(_07701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15798_ (.A1(_06798_),
    .A2(_07659_),
    .B(_07701_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15799_ (.A1(_06806_),
    .A2(_07698_),
    .ZN(_07702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15800_ (.I(_07649_),
    .Z(_07703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15801_ (.I(_07663_),
    .Z(_07704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15802_ (.A1(\filters.low[18] ),
    .A2(_07703_),
    .B(_07704_),
    .ZN(_07705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15803_ (.A1(_07702_),
    .A2(_07705_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15804_ (.A1(_06814_),
    .A2(_07698_),
    .ZN(_07706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15805_ (.A1(\filters.low[19] ),
    .A2(_07703_),
    .B(_07704_),
    .ZN(_07707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15806_ (.A1(_07706_),
    .A2(_07707_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15807_ (.A1(_06824_),
    .A2(_07698_),
    .ZN(_07708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15808_ (.A1(\filters.low[20] ),
    .A2(_07703_),
    .B(_07704_),
    .ZN(_07709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15809_ (.A1(_07708_),
    .A2(_07709_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15810_ (.I(_07682_),
    .Z(_07710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15811_ (.A1(_06834_),
    .A2(_07710_),
    .ZN(_07711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15812_ (.A1(_07350_),
    .A2(_07703_),
    .B(_07704_),
    .ZN(_07712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15813_ (.A1(_07711_),
    .A2(_07712_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15814_ (.A1(_06842_),
    .A2(_07710_),
    .ZN(_07713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15815_ (.I(_07649_),
    .Z(_07714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15816_ (.I(_01761_),
    .Z(_07715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15817_ (.I(_07715_),
    .Z(_07716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15818_ (.A1(\filters.low[22] ),
    .A2(_07714_),
    .B(_07716_),
    .ZN(_07717_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15819_ (.A1(_07713_),
    .A2(_07717_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15820_ (.I(_07655_),
    .Z(_07718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15821_ (.I(_07682_),
    .Z(_07719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15822_ (.A1(_06852_),
    .A2(_07719_),
    .ZN(_07720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15823_ (.A1(_06846_),
    .A2(_07718_),
    .B(_07720_),
    .C(_07219_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15824_ (.A1(_07381_),
    .A2(_07650_),
    .B(_07688_),
    .ZN(_07721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15825_ (.A1(_06865_),
    .A2(_07659_),
    .B(_07721_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15826_ (.A1(_06872_),
    .A2(_07710_),
    .ZN(_07722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15827_ (.A1(_07391_),
    .A2(_07714_),
    .B(_07716_),
    .ZN(_07723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15828_ (.A1(_07722_),
    .A2(_07723_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15829_ (.A1(_06883_),
    .A2(_07710_),
    .ZN(_07724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15830_ (.A1(_07401_),
    .A2(_07714_),
    .B(_07716_),
    .ZN(_07725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15831_ (.A1(_07724_),
    .A2(_07725_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15832_ (.A1(_06891_),
    .A2(_07719_),
    .ZN(_07726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15833_ (.A1(_07413_),
    .A2(_07714_),
    .B(_07716_),
    .ZN(_07727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15834_ (.A1(_07726_),
    .A2(_07727_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15835_ (.A1(_06903_),
    .A2(_07719_),
    .ZN(_07728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15836_ (.I(_02355_),
    .Z(_07729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15837_ (.A1(_06899_),
    .A2(_07718_),
    .B(_07728_),
    .C(_07729_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15838_ (.A1(_06912_),
    .A2(_07719_),
    .ZN(_07730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15839_ (.A1(_06906_),
    .A2(_07718_),
    .B(_07730_),
    .C(_07729_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15840_ (.A1(_06922_),
    .A2(_07655_),
    .ZN(_07731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15841_ (.A1(_06916_),
    .A2(_07718_),
    .B(_07731_),
    .C(_07729_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15842_ (.A1(\filters.low[31] ),
    .A2(_07650_),
    .B(_07688_),
    .ZN(_07732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15843_ (.A1(_06929_),
    .A2(_07659_),
    .B(_07732_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15844_ (.I(_03761_),
    .Z(_07733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15845_ (.A1(_07733_),
    .A2(_07647_),
    .ZN(_07734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15846_ (.A1(_04242_),
    .A2(_04186_),
    .B(_07734_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15847_ (.A1(_03216_),
    .A2(_03218_),
    .A3(_03759_),
    .ZN(_07735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15848_ (.A1(_07733_),
    .A2(_07735_),
    .ZN(_07736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15849_ (.A1(_03196_),
    .A2(_07647_),
    .B(_07736_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15850_ (.A1(_07461_),
    .A2(_07735_),
    .Z(_07737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15851_ (.A1(_07617_),
    .A2(_07737_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15852_ (.A1(\spi_dac_i.counter[4] ),
    .A2(\spi_dac_i.counter[3] ),
    .Z(_07738_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15853_ (.A1(\spi_dac_i.counter[0] ),
    .A2(_07738_),
    .Z(_07739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15854_ (.I(_07739_),
    .Z(_07740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15855_ (.I(\spi_dac_i.counter[0] ),
    .Z(_07741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15856_ (.I(_07738_),
    .Z(_07742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15857_ (.I(_07742_),
    .Z(_07743_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15858_ (.A1(_07741_),
    .A2(_04809_),
    .A3(_07743_),
    .ZN(_07744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15859_ (.I(_07566_),
    .Z(_07745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15860_ (.A1(_07740_),
    .A2(_07744_),
    .B(_07745_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15861_ (.I(\spi_dac_i.counter[3] ),
    .Z(_07746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15862_ (.A1(\spi_dac_i.counter[4] ),
    .A2(_07746_),
    .ZN(_07747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15863_ (.I(_07747_),
    .Z(_07748_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15864_ (.A1(\spi_dac_i.counter[0] ),
    .A2(_07748_),
    .Z(_07749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15865_ (.I(_07749_),
    .Z(_07750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15866_ (.I(_07739_),
    .Z(_07751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15867_ (.A1(_04809_),
    .A2(_07742_),
    .ZN(_07752_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15868_ (.A1(\spi_dac_i.counter[1] ),
    .A2(_07751_),
    .A3(_07752_),
    .ZN(_07753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15869_ (.A1(\spi_dac_i.counter[1] ),
    .A2(_07750_),
    .B(_07753_),
    .ZN(_07754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15870_ (.A1(_07617_),
    .A2(_07754_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _15871_ (.A1(\spi_dac_i.counter[2] ),
    .A2(\spi_dac_i.counter[1] ),
    .A3(_07741_),
    .Z(_07755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15872_ (.A1(\spi_dac_i.counter[1] ),
    .A2(_07741_),
    .B(\spi_dac_i.counter[2] ),
    .ZN(_07756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15873_ (.I(\spi_dac_i.counter[2] ),
    .ZN(_07757_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _15874_ (.A1(_07742_),
    .A2(_07755_),
    .A3(_07756_),
    .B1(_07752_),
    .B2(_07757_),
    .ZN(_07758_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15875_ (.A1(_07733_),
    .A2(_07758_),
    .Z(_07759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15876_ (.I(_07759_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15877_ (.A1(\spi_dac_i.counter[4] ),
    .A2(_07755_),
    .B(_07746_),
    .ZN(_07760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15878_ (.A1(_07746_),
    .A2(_07755_),
    .B(_07760_),
    .ZN(_07761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15879_ (.A1(_07752_),
    .A2(_07761_),
    .B(_07745_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15880_ (.I(_07738_),
    .Z(_07762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15881_ (.I(_07762_),
    .Z(_07763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15882_ (.I(_07763_),
    .Z(_07764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15883_ (.A1(_07746_),
    .A2(_07755_),
    .B(\spi_dac_i.counter[4] ),
    .ZN(_07765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _15884_ (.A1(_04198_),
    .A2(_07764_),
    .B(_07765_),
    .C(_07729_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15885_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.in ),
    .ZN(_07766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15886_ (.I(_07766_),
    .Z(_07767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15887_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ),
    .A2(_07767_),
    .ZN(_07768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _15888_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ),
    .A2(_07767_),
    .ZN(_07769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15889_ (.I(_07769_),
    .Z(_07770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15890_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ),
    .A2(_07766_),
    .ZN(_07771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15891_ (.I(_07771_),
    .Z(_07772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15892_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ),
    .A2(_07770_),
    .ZN(_07773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15893_ (.A1(_07770_),
    .A2(_07772_),
    .B(_07773_),
    .ZN(_07774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15894_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ),
    .A2(_07767_),
    .ZN(_07775_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15895_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ),
    .ZN(_07776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15896_ (.A1(_07776_),
    .A2(\tt_um_rejunity_sn76489.chan[2].attenuation.in ),
    .ZN(_07777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15897_ (.I(_07777_),
    .Z(_07778_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15898_ (.A1(_07778_),
    .A2(_07772_),
    .Z(_07779_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15899_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ),
    .ZN(_07780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15900_ (.A1(_07780_),
    .A2(_02349_),
    .ZN(_07781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15901_ (.I(_07781_),
    .Z(_07782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15902_ (.A1(_07775_),
    .A2(_07779_),
    .B(_07782_),
    .ZN(_07783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15903_ (.I(_07783_),
    .ZN(_07784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15904_ (.A1(_07768_),
    .A2(_07774_),
    .B(_07784_),
    .ZN(_07785_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15905_ (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.in ),
    .ZN(_07786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15906_ (.I(_07786_),
    .Z(_07787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15907_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ),
    .A2(_07787_),
    .ZN(_07788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15908_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ),
    .A2(_07786_),
    .ZN(_07789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15909_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ),
    .A2(_07787_),
    .ZN(_07790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15910_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ),
    .A2(_07789_),
    .ZN(_07791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15911_ (.A1(_07789_),
    .A2(_07790_),
    .B(_07791_),
    .ZN(_07792_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15912_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ),
    .A2(_07786_),
    .Z(_07793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15913_ (.I(_07793_),
    .Z(_07794_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15914_ (.I(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ),
    .ZN(_07795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15915_ (.A1(_07795_),
    .A2(\tt_um_rejunity_sn76489.chan[1].attenuation.in ),
    .ZN(_07796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15916_ (.A1(_07794_),
    .A2(_07796_),
    .ZN(_07797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15917_ (.I(_07789_),
    .Z(_07798_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15918_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ),
    .A2(_07787_),
    .Z(_07799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15919_ (.A1(_07798_),
    .A2(_07790_),
    .B(_07799_),
    .ZN(_07800_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15920_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ),
    .A2(_07787_),
    .Z(_07801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15921_ (.A1(_07797_),
    .A2(_07800_),
    .B(_07801_),
    .ZN(_07802_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15922_ (.I(_07802_),
    .ZN(_07803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15923_ (.A1(_07788_),
    .A2(_07792_),
    .B(_07803_),
    .ZN(_07804_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _15924_ (.I(\tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ),
    .ZN(_07805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15925_ (.A1(_07805_),
    .A2(\tt_um_rejunity_sn76489.chan[0].attenuation.in ),
    .ZN(_07806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15926_ (.I(_07806_),
    .Z(_07807_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15927_ (.I(\tt_um_rejunity_sn76489.chan[0].attenuation.in ),
    .ZN(_07808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15928_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ),
    .A2(_07808_),
    .ZN(_07809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15929_ (.A1(_07807_),
    .A2(_07809_),
    .ZN(_07810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15930_ (.I(_07808_),
    .Z(_07811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15931_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ),
    .A2(_07811_),
    .ZN(_07812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15932_ (.I(_07812_),
    .Z(_07813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15933_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ),
    .A2(_07811_),
    .ZN(_07814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15934_ (.I(_07814_),
    .Z(_07815_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _15935_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ),
    .A2(_07811_),
    .Z(_07816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15936_ (.A1(_07813_),
    .A2(_07815_),
    .B(_07816_),
    .ZN(_07817_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15937_ (.I(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ),
    .ZN(_07818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15938_ (.I(\tt_um_rejunity_sn76489.chan[0].attenuation.in ),
    .Z(_07819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15939_ (.A1(_07818_),
    .A2(_07819_),
    .ZN(_07820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15940_ (.A1(_07806_),
    .A2(_07820_),
    .ZN(_07821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15941_ (.I(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ),
    .Z(_07822_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _15942_ (.A1(_07805_),
    .A2(_07818_),
    .B(_07822_),
    .C(_07819_),
    .ZN(_07823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15943_ (.A1(_07821_),
    .A2(_07823_),
    .B(_07816_),
    .ZN(_07824_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15944_ (.I(_07824_),
    .ZN(_07825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _15945_ (.A1(_07810_),
    .A2(_07817_),
    .B(_07825_),
    .ZN(_07826_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _15946_ (.A1(_07804_),
    .A2(_07826_),
    .ZN(_07827_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15947_ (.I(_07827_),
    .ZN(_07828_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15948_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.in ),
    .ZN(_07829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15949_ (.I(_07829_),
    .Z(_07830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15950_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ),
    .A2(_07830_),
    .ZN(_07831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15951_ (.I(_07831_),
    .Z(_07832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15952_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ),
    .A2(_07829_),
    .ZN(_07833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15953_ (.I(_07833_),
    .Z(_07834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15954_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ),
    .A2(_07830_),
    .ZN(_07835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15955_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ),
    .A2(_07833_),
    .ZN(_07836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _15956_ (.A1(_07834_),
    .A2(_07835_),
    .B(_07836_),
    .ZN(_07837_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _15957_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ),
    .ZN(_07838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15958_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.in ),
    .Z(_07839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15959_ (.A1(_07838_),
    .A2(_07839_),
    .ZN(_07840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15960_ (.I(_07840_),
    .Z(_07841_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15961_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ),
    .ZN(_07842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15962_ (.A1(_07842_),
    .A2(_07839_),
    .ZN(_07843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15963_ (.I(_07843_),
    .Z(_07844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15964_ (.A1(_07841_),
    .A2(_07844_),
    .ZN(_07845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15965_ (.I(_07834_),
    .Z(_07846_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _15966_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ),
    .ZN(_07847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _15967_ (.A1(_07847_),
    .A2(\tt_um_rejunity_sn76489.chan[3].attenuation.in ),
    .ZN(_07848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _15968_ (.A1(_07846_),
    .A2(_07835_),
    .B(_07848_),
    .ZN(_07849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15969_ (.A1(_07845_),
    .A2(_07849_),
    .ZN(_07850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15970_ (.A1(_07831_),
    .A2(_07850_),
    .ZN(_07851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _15971_ (.A1(_07832_),
    .A2(_07837_),
    .B(_07851_),
    .ZN(_07852_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _15972_ (.A1(_07828_),
    .A2(_07852_),
    .Z(_07853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15973_ (.A1(_07785_),
    .A2(_07853_),
    .ZN(_07854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _15974_ (.I(_07748_),
    .Z(_07855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15975_ (.A1(_07785_),
    .A2(_07853_),
    .ZN(_07856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15976_ (.A1(_07855_),
    .A2(_07856_),
    .ZN(_07857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _15977_ (.A1(\spi_dac_i.spi_dat_buff_1[0] ),
    .A2(_07750_),
    .B1(_07854_),
    .B2(_07857_),
    .ZN(_07858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15978_ (.A1(_07617_),
    .A2(_07858_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15979_ (.I(_07743_),
    .Z(_07859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15980_ (.A1(_07828_),
    .A2(_07852_),
    .ZN(_07860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15981_ (.A1(_07860_),
    .A2(_07854_),
    .ZN(_07861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _15982_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ),
    .Z(_07862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15983_ (.A1(_07768_),
    .A2(_07773_),
    .ZN(_07863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15984_ (.A1(_07778_),
    .A2(_07775_),
    .ZN(_07864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15985_ (.A1(_07782_),
    .A2(_07864_),
    .ZN(_07865_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _15986_ (.A1(_07862_),
    .A2(_07863_),
    .B1(_07865_),
    .B2(_07774_),
    .ZN(_07866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15987_ (.A1(_07834_),
    .A2(_07848_),
    .ZN(_07867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15988_ (.A1(_07831_),
    .A2(_07836_),
    .ZN(_07868_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _15989_ (.A1(_07831_),
    .A2(_07837_),
    .A3(_07867_),
    .B1(_07868_),
    .B2(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ),
    .ZN(_07869_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _15990_ (.A1(_07804_),
    .A2(_07826_),
    .Z(_07870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15991_ (.A1(_07822_),
    .A2(_07812_),
    .ZN(_07871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15992_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ),
    .A2(_07809_),
    .ZN(_07872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15993_ (.A1(_07816_),
    .A2(_07807_),
    .A3(_07872_),
    .ZN(_07873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _15994_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ),
    .A2(_07811_),
    .ZN(_07874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15995_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ),
    .A2(_07874_),
    .ZN(_07875_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _15996_ (.A1(_07871_),
    .A2(_07873_),
    .A3(_07875_),
    .ZN(_07876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15997_ (.A1(_07788_),
    .A2(_07791_),
    .ZN(_07877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _15998_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ),
    .A2(_07786_),
    .ZN(_07878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _15999_ (.A1(_07793_),
    .A2(_07878_),
    .ZN(_07879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16000_ (.A1(_07801_),
    .A2(_07879_),
    .ZN(_07880_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _16001_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ),
    .A2(_07877_),
    .B1(_07880_),
    .B2(_07792_),
    .ZN(_07881_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16002_ (.A1(_07876_),
    .A2(_07881_),
    .Z(_07882_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16003_ (.I(_07882_),
    .ZN(_07883_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16004_ (.A1(_07870_),
    .A2(_07883_),
    .Z(_07884_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16005_ (.A1(_07869_),
    .A2(_07884_),
    .Z(_07885_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16006_ (.A1(_07866_),
    .A2(_07885_),
    .ZN(_07886_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16007_ (.A1(_07861_),
    .A2(_07886_),
    .Z(_07887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16008_ (.I(_07751_),
    .Z(_07888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16009_ (.A1(\spi_dac_i.counter[0] ),
    .A2(_07747_),
    .ZN(_07889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16010_ (.I(_07889_),
    .Z(_07890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16011_ (.I(_07890_),
    .Z(_07891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16012_ (.I(_03508_),
    .Z(_07892_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16013_ (.A1(\spi_dac_i.spi_dat_buff_1[0] ),
    .A2(_07888_),
    .B1(_07891_),
    .B2(\spi_dac_i.spi_dat_buff_1[1] ),
    .C(_07892_),
    .ZN(_07893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16014_ (.A1(_07859_),
    .A2(_07887_),
    .B(_07893_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16015_ (.A1(_07860_),
    .A2(_07854_),
    .B(_07886_),
    .ZN(_07894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16016_ (.A1(_07771_),
    .A2(_07775_),
    .ZN(_07895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16017_ (.I(_07895_),
    .Z(_07896_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _16018_ (.A1(_07862_),
    .A2(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ),
    .A3(_07767_),
    .ZN(_07897_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _16019_ (.A1(_07769_),
    .A2(_07895_),
    .A3(_07897_),
    .ZN(_07898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16020_ (.A1(_07777_),
    .A2(_07772_),
    .ZN(_07899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16021_ (.A1(_07768_),
    .A2(_07899_),
    .ZN(_07900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _16022_ (.A1(_07769_),
    .A2(_07896_),
    .B(_07898_),
    .C(_07900_),
    .ZN(_07901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16023_ (.A1(_07809_),
    .A2(_07815_),
    .ZN(_07902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16024_ (.A1(_07809_),
    .A2(_07814_),
    .ZN(_07903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16025_ (.A1(_07813_),
    .A2(_07903_),
    .ZN(_07904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16026_ (.A1(_07902_),
    .A2(_07904_),
    .ZN(_07905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16027_ (.A1(_07820_),
    .A2(_07815_),
    .ZN(_07906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16028_ (.A1(_07812_),
    .A2(_07820_),
    .ZN(_07907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16029_ (.A1(_07874_),
    .A2(_07907_),
    .ZN(_07908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16030_ (.A1(_07906_),
    .A2(_07908_),
    .ZN(_07909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16031_ (.A1(_07905_),
    .A2(_07909_),
    .ZN(_07910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16032_ (.I(_07796_),
    .Z(_07911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16033_ (.A1(_07911_),
    .A2(_07799_),
    .ZN(_07912_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16034_ (.A1(_07790_),
    .A2(_07878_),
    .Z(_07913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16035_ (.A1(_07798_),
    .A2(_07911_),
    .B(_07788_),
    .ZN(_07914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16036_ (.A1(_07794_),
    .A2(_07913_),
    .B(_07914_),
    .ZN(_07915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16037_ (.A1(_07794_),
    .A2(_07912_),
    .B(_07915_),
    .ZN(_07916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16038_ (.A1(_07910_),
    .A2(_07916_),
    .ZN(_07917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16039_ (.I(_07917_),
    .ZN(_07918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16040_ (.A1(_07910_),
    .A2(_07916_),
    .ZN(_07919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16041_ (.A1(_07918_),
    .A2(_07919_),
    .ZN(_07920_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _16042_ (.A1(_07871_),
    .A2(_07873_),
    .A3(_07875_),
    .A4(_07881_),
    .ZN(_07921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16043_ (.A1(_07870_),
    .A2(_07883_),
    .ZN(_07922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16044_ (.A1(_07921_),
    .A2(_07922_),
    .ZN(_07923_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16045_ (.A1(_07920_),
    .A2(_07923_),
    .ZN(_07924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16046_ (.A1(_07843_),
    .A2(_07848_),
    .ZN(_07925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16047_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ),
    .A2(_07830_),
    .ZN(_07926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16048_ (.A1(_07835_),
    .A2(_07926_),
    .ZN(_07927_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16049_ (.A1(_07925_),
    .A2(_07927_),
    .Z(_07928_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16050_ (.A1(_07840_),
    .A2(_07928_),
    .Z(_07929_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _16051_ (.I(\tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ),
    .ZN(_07930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16052_ (.A1(_07930_),
    .A2(_07839_),
    .ZN(_07931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16053_ (.A1(_07834_),
    .A2(_07843_),
    .ZN(_07932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16054_ (.A1(_07931_),
    .A2(_07932_),
    .ZN(_07933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16055_ (.A1(_07841_),
    .A2(_07925_),
    .B(_07933_),
    .ZN(_07934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16056_ (.A1(_07929_),
    .A2(_07934_),
    .ZN(_07935_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _16057_ (.A1(_07901_),
    .A2(_07924_),
    .A3(_07935_),
    .Z(_07936_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16058_ (.I(_07936_),
    .ZN(_07937_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16059_ (.A1(_07869_),
    .A2(_07884_),
    .Z(_07938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16060_ (.A1(_07866_),
    .A2(_07885_),
    .B(_07938_),
    .ZN(_07939_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16061_ (.A1(_07937_),
    .A2(_07939_),
    .Z(_07940_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16062_ (.A1(_07894_),
    .A2(_07940_),
    .ZN(_07941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16063_ (.I(_07889_),
    .Z(_07942_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16064_ (.A1(\spi_dac_i.spi_dat_buff_1[1] ),
    .A2(_07888_),
    .B1(_07942_),
    .B2(\spi_dac_i.spi_dat_buff_1[2] ),
    .C(_07892_),
    .ZN(_07943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16065_ (.A1(_07859_),
    .A2(_07941_),
    .B(_07943_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16066_ (.I(_07616_),
    .Z(_07944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16067_ (.I(_07890_),
    .Z(_07945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16068_ (.A1(_07894_),
    .A2(_07940_),
    .ZN(_07946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16069_ (.A1(_07937_),
    .A2(_07939_),
    .B(_07946_),
    .ZN(_07947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16070_ (.A1(_07781_),
    .A2(_07896_),
    .ZN(_07948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16071_ (.A1(_07862_),
    .A2(_07775_),
    .ZN(_07949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _16072_ (.A1(\tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ),
    .A2(_07948_),
    .B1(_07949_),
    .B2(_07781_),
    .C(_07899_),
    .ZN(_07950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16073_ (.I(_07874_),
    .Z(_07951_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _16074_ (.A1(_07805_),
    .A2(_07951_),
    .A3(_07906_),
    .B1(_07908_),
    .B2(_07904_),
    .ZN(_07952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16075_ (.A1(_07798_),
    .A2(_07911_),
    .ZN(_07953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16076_ (.I(_07788_),
    .Z(_07954_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16077_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ),
    .A2(_07954_),
    .A3(_07912_),
    .ZN(_07955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16078_ (.A1(_07795_),
    .A2(_07799_),
    .B(_07801_),
    .ZN(_07956_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _16079_ (.A1(_07953_),
    .A2(_07955_),
    .A3(_07956_),
    .ZN(_07957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16080_ (.A1(_07917_),
    .A2(_07923_),
    .B(_07919_),
    .ZN(_07958_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _16081_ (.A1(_07952_),
    .A2(_07957_),
    .A3(_07958_),
    .Z(_07959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16082_ (.A1(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ),
    .A2(_07926_),
    .ZN(_07960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16083_ (.I(_07931_),
    .Z(_07961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _16084_ (.A1(_07844_),
    .A2(_07848_),
    .B(_07838_),
    .C(_07931_),
    .ZN(_07962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _16085_ (.A1(_07846_),
    .A2(_07844_),
    .B1(_07960_),
    .B2(_07961_),
    .C(_07962_),
    .ZN(_07963_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _16086_ (.A1(_07950_),
    .A2(_07959_),
    .A3(_07963_),
    .ZN(_07964_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16087_ (.A1(_07924_),
    .A2(_07935_),
    .Z(_07965_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16088_ (.A1(_07924_),
    .A2(_07935_),
    .Z(_07966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16089_ (.A1(_07901_),
    .A2(_07965_),
    .B(_07966_),
    .ZN(_07967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16090_ (.A1(_07964_),
    .A2(_07967_),
    .Z(_07968_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16091_ (.A1(_07947_),
    .A2(_07968_),
    .Z(_07969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16092_ (.A1(_07947_),
    .A2(_07968_),
    .B(_07742_),
    .ZN(_07970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16093_ (.A1(\spi_dac_i.spi_dat_buff_1[2] ),
    .A2(_07748_),
    .ZN(_07971_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16094_ (.A1(_07969_),
    .A2(_07970_),
    .B(_07971_),
    .C(_07890_),
    .ZN(_07972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16095_ (.A1(\spi_dac_i.spi_dat_buff_1[3] ),
    .A2(_07945_),
    .B(_07972_),
    .ZN(_07973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16096_ (.A1(_07944_),
    .A2(_07973_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16097_ (.A1(_07964_),
    .A2(_07967_),
    .ZN(_07974_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16098_ (.A1(_07974_),
    .A2(_07969_),
    .Z(_07975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16099_ (.I(_07897_),
    .Z(_07976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16100_ (.A1(_07782_),
    .A2(_07976_),
    .B(_07783_),
    .ZN(_07977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16101_ (.A1(_07832_),
    .A2(_07927_),
    .ZN(_07978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16102_ (.A1(_07832_),
    .A2(_07850_),
    .B(_07978_),
    .ZN(_07979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16103_ (.A1(_07951_),
    .A2(_07902_),
    .B(_07825_),
    .ZN(_07980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16104_ (.I(_07801_),
    .Z(_07981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16105_ (.A1(_07911_),
    .A2(_07799_),
    .ZN(_07982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16106_ (.A1(_07981_),
    .A2(_07982_),
    .B(_07802_),
    .ZN(_07983_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16107_ (.A1(_07980_),
    .A2(_07983_),
    .ZN(_07984_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16108_ (.I(_07952_),
    .ZN(_07985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16109_ (.A1(_07985_),
    .A2(_07957_),
    .ZN(_07986_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16110_ (.A1(_07917_),
    .A2(_07923_),
    .A3(_07986_),
    .ZN(_07987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16111_ (.A1(_07985_),
    .A2(_07957_),
    .B(_07987_),
    .ZN(_07988_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16112_ (.A1(_07984_),
    .A2(_07988_),
    .ZN(_07989_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _16113_ (.A1(_07977_),
    .A2(_07979_),
    .A3(_07989_),
    .Z(_07990_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16114_ (.A1(_07959_),
    .A2(_07963_),
    .Z(_07991_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16115_ (.A1(_07959_),
    .A2(_07963_),
    .Z(_07992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16116_ (.A1(_07950_),
    .A2(_07991_),
    .B(_07992_),
    .ZN(_07993_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _16117_ (.A1(_07975_),
    .A2(_07990_),
    .A3(_07993_),
    .ZN(_07994_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16118_ (.A1(\spi_dac_i.spi_dat_buff_1[3] ),
    .A2(_07888_),
    .B1(_07942_),
    .B2(\spi_dac_i.spi_dat_buff_1[4] ),
    .C(_07892_),
    .ZN(_07995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16119_ (.A1(_07859_),
    .A2(_07994_),
    .B(_07995_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16120_ (.A1(_07990_),
    .A2(_07993_),
    .ZN(_07996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16121_ (.A1(_07990_),
    .A2(_07993_),
    .ZN(_07997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16122_ (.A1(_07975_),
    .A2(_07996_),
    .B(_07997_),
    .ZN(_07998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16123_ (.I(_07977_),
    .ZN(_07999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16124_ (.A1(_07979_),
    .A2(_07989_),
    .ZN(_08000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16125_ (.A1(_07979_),
    .A2(_07989_),
    .ZN(_08001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16126_ (.A1(_07999_),
    .A2(_08000_),
    .B(_08001_),
    .ZN(_08002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16127_ (.A1(_07770_),
    .A2(_07772_),
    .ZN(_08003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16128_ (.I(_07768_),
    .Z(_08004_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16129_ (.A1(_08004_),
    .A2(_07896_),
    .A3(_07976_),
    .ZN(_08005_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16130_ (.A1(_08003_),
    .A2(_08005_),
    .ZN(_08006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16131_ (.A1(_07961_),
    .A2(_07928_),
    .ZN(_08007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16132_ (.A1(_07845_),
    .A2(_08007_),
    .Z(_08008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16133_ (.I(_07816_),
    .Z(_08009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16134_ (.A1(_08009_),
    .A2(_07902_),
    .ZN(_08010_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16135_ (.A1(_07903_),
    .A2(_08010_),
    .Z(_08011_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16136_ (.A1(_07821_),
    .A2(_08011_),
    .ZN(_08012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16137_ (.A1(_07981_),
    .A2(_07913_),
    .ZN(_08013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16138_ (.A1(_07797_),
    .A2(_08013_),
    .ZN(_08014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16139_ (.A1(_08012_),
    .A2(_08014_),
    .ZN(_08015_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16140_ (.A1(_08012_),
    .A2(_08014_),
    .Z(_08016_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16141_ (.A1(_08015_),
    .A2(_08016_),
    .Z(_08017_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _16142_ (.A1(_07981_),
    .A2(_07982_),
    .B(_07980_),
    .C(_07802_),
    .ZN(_08018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16143_ (.A1(_07984_),
    .A2(_07988_),
    .ZN(_08019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16144_ (.A1(_08018_),
    .A2(_08019_),
    .ZN(_08020_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16145_ (.A1(_08017_),
    .A2(_08020_),
    .ZN(_08021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16146_ (.A1(_08008_),
    .A2(_08021_),
    .Z(_08022_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16147_ (.A1(_08006_),
    .A2(_08022_),
    .ZN(_08023_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _16148_ (.A1(_07998_),
    .A2(_08002_),
    .A3(_08023_),
    .Z(_08024_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16149_ (.A1(\spi_dac_i.spi_dat_buff_1[4] ),
    .A2(_07888_),
    .B1(_07942_),
    .B2(\spi_dac_i.spi_dat_buff_1[5] ),
    .C(_07892_),
    .ZN(_08025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16150_ (.A1(_07764_),
    .A2(_08024_),
    .B(_08025_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16151_ (.A1(_08002_),
    .A2(_08023_),
    .Z(_08026_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16152_ (.A1(_08002_),
    .A2(_08023_),
    .Z(_08027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16153_ (.A1(_07998_),
    .A2(_08026_),
    .B(_08027_),
    .ZN(_08028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16154_ (.A1(_07778_),
    .A2(_07976_),
    .B(_07864_),
    .ZN(_08029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16155_ (.A1(_07778_),
    .A2(_07976_),
    .ZN(_08030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16156_ (.A1(_08004_),
    .A2(_08029_),
    .B1(_08030_),
    .B2(_07900_),
    .ZN(_08031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16157_ (.A1(_07846_),
    .A2(_07927_),
    .B(_07867_),
    .ZN(_08032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16158_ (.A1(_07846_),
    .A2(_07927_),
    .ZN(_08033_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _16159_ (.A1(_07961_),
    .A2(_08032_),
    .B1(_08033_),
    .B2(_07933_),
    .ZN(_08034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16160_ (.I(_07794_),
    .Z(_08035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16161_ (.A1(_08035_),
    .A2(_07982_),
    .B(_07879_),
    .ZN(_08036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16162_ (.A1(_08035_),
    .A2(_07982_),
    .ZN(_08037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _16163_ (.A1(_07954_),
    .A2(_08036_),
    .B1(_08037_),
    .B2(_07914_),
    .ZN(_08038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16164_ (.A1(_07822_),
    .A2(_07807_),
    .B1(_07821_),
    .B2(_07815_),
    .ZN(_08039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16165_ (.A1(_07813_),
    .A2(_07902_),
    .B(_07907_),
    .ZN(_08040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16166_ (.A1(_08009_),
    .A2(_08040_),
    .ZN(_08041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16167_ (.A1(_08009_),
    .A2(_08039_),
    .B(_08041_),
    .ZN(_08042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16168_ (.A1(_08017_),
    .A2(_08020_),
    .ZN(_08043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16169_ (.A1(_08015_),
    .A2(_08043_),
    .ZN(_08044_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _16170_ (.A1(_08038_),
    .A2(_08042_),
    .A3(_08044_),
    .ZN(_08045_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16171_ (.A1(_08034_),
    .A2(_08045_),
    .ZN(_08046_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16172_ (.A1(_08031_),
    .A2(_08046_),
    .ZN(_08047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16173_ (.A1(_08006_),
    .A2(_08022_),
    .ZN(_08048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16174_ (.A1(_08008_),
    .A2(_08021_),
    .B(_08048_),
    .ZN(_08049_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _16175_ (.A1(_08028_),
    .A2(_08047_),
    .A3(_08049_),
    .ZN(_08050_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16176_ (.A1(\spi_dac_i.spi_dat_buff_1[5] ),
    .A2(_07751_),
    .B1(_07942_),
    .B2(\spi_dac_i.spi_dat_buff_1[6] ),
    .C(_03761_),
    .ZN(_08051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16177_ (.A1(_07764_),
    .A2(_08050_),
    .B(_08051_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16178_ (.A1(_08047_),
    .A2(_08049_),
    .Z(_08052_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16179_ (.A1(_08047_),
    .A2(_08049_),
    .Z(_08053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16180_ (.A1(_08028_),
    .A2(_08052_),
    .B(_08053_),
    .ZN(_08054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _16181_ (.A1(_08004_),
    .A2(_08029_),
    .B1(_08030_),
    .B2(_07900_),
    .C(_08046_),
    .ZN(_08055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16182_ (.I(_08055_),
    .ZN(_08056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16183_ (.A1(_08034_),
    .A2(_08045_),
    .B(_08056_),
    .ZN(_08057_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _16184_ (.A1(_07780_),
    .A2(_08003_),
    .B1(_07863_),
    .B2(_07898_),
    .ZN(_08058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16185_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ),
    .A2(_07821_),
    .ZN(_08059_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16186_ (.A1(_07951_),
    .A2(_07871_),
    .A3(_07905_),
    .ZN(_08060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16187_ (.A1(_08035_),
    .A2(_07913_),
    .B(_07877_),
    .ZN(_08061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16188_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ),
    .A2(_07797_),
    .B(_08061_),
    .ZN(_08062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16189_ (.A1(_08059_),
    .A2(_08060_),
    .B(_08062_),
    .ZN(_08063_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16190_ (.A1(_08062_),
    .A2(_08059_),
    .A3(_08060_),
    .Z(_08064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16191_ (.A1(_08063_),
    .A2(_08064_),
    .ZN(_08065_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16192_ (.A1(_08038_),
    .A2(_08042_),
    .Z(_08066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16193_ (.A1(_08038_),
    .A2(_08042_),
    .ZN(_08067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16194_ (.I(_08067_),
    .ZN(_08068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16195_ (.A1(_08066_),
    .A2(_08044_),
    .B(_08068_),
    .ZN(_08069_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16196_ (.A1(_08065_),
    .A2(_08069_),
    .ZN(_08070_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _16197_ (.A1(_07930_),
    .A2(_07841_),
    .A3(_07844_),
    .B1(_07868_),
    .B2(_07929_),
    .ZN(_08071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16198_ (.A1(_08070_),
    .A2(_08071_),
    .Z(_08072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16199_ (.A1(_08058_),
    .A2(_08072_),
    .Z(_08073_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _16200_ (.A1(_08054_),
    .A2(_08057_),
    .A3(_08073_),
    .Z(_08074_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16201_ (.A1(\spi_dac_i.spi_dat_buff_1[6] ),
    .A2(_07751_),
    .B1(_07890_),
    .B2(\spi_dac_i.spi_dat_buff_1[7] ),
    .C(_03761_),
    .ZN(_08075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16202_ (.A1(_07764_),
    .A2(_08074_),
    .B(_08075_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16203_ (.A1(_08057_),
    .A2(_08073_),
    .ZN(_08076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16204_ (.A1(_08057_),
    .A2(_08073_),
    .ZN(_08077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16205_ (.A1(_08054_),
    .A2(_08076_),
    .B(_08077_),
    .ZN(_08078_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _16206_ (.A1(_07782_),
    .A2(_07896_),
    .A3(_07899_),
    .ZN(_08079_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _16207_ (.A1(_07832_),
    .A2(_07925_),
    .A3(_07932_),
    .ZN(_08080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16208_ (.I(_08016_),
    .ZN(_08081_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _16209_ (.A1(_08018_),
    .A2(_08081_),
    .B(_08067_),
    .C(_08015_),
    .ZN(_08082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16210_ (.A1(_08038_),
    .A2(_08042_),
    .ZN(_08083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16211_ (.A1(_08083_),
    .A2(_08064_),
    .ZN(_08084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16212_ (.A1(_08082_),
    .A2(_08084_),
    .B(_08063_),
    .ZN(_08085_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _16213_ (.A1(_07954_),
    .A2(_07912_),
    .A3(_07953_),
    .ZN(_08086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16214_ (.A1(_07903_),
    .A2(_07908_),
    .ZN(_08087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16215_ (.A1(_08086_),
    .A2(_08087_),
    .Z(_08088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16216_ (.A1(_08085_),
    .A2(_08088_),
    .ZN(_08089_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _16217_ (.A1(_08079_),
    .A2(_08080_),
    .A3(_08089_),
    .ZN(_08090_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16218_ (.A1(_08070_),
    .A2(_08071_),
    .Z(_08091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16219_ (.A1(_08058_),
    .A2(_08072_),
    .B(_08091_),
    .ZN(_08092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16220_ (.A1(_08090_),
    .A2(_08092_),
    .Z(_08093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16221_ (.A1(_08078_),
    .A2(_08093_),
    .Z(_08094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16222_ (.A1(_07855_),
    .A2(_08094_),
    .ZN(_08095_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _16223_ (.A1(\spi_dac_i.spi_dat_buff_1[7] ),
    .A2(_07740_),
    .B1(_07891_),
    .B2(\spi_dac_i.spi_dat_buff_1[8] ),
    .C(_03509_),
    .ZN(_08096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16224_ (.A1(_08095_),
    .A2(_08096_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16225_ (.A1(_08078_),
    .A2(_08093_),
    .ZN(_08097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16226_ (.A1(_08090_),
    .A2(_08092_),
    .B(_08097_),
    .ZN(_08098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16227_ (.A1(_08004_),
    .A2(_07770_),
    .ZN(_08099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16228_ (.A1(_07961_),
    .A2(_07841_),
    .ZN(_08100_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16229_ (.A1(_07903_),
    .A2(_07908_),
    .A3(_08086_),
    .ZN(_08101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16230_ (.A1(_08085_),
    .A2(_08088_),
    .ZN(_08102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16231_ (.A1(_08101_),
    .A2(_08102_),
    .ZN(_08103_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _16232_ (.A1(_07954_),
    .A2(_07798_),
    .A3(_07951_),
    .A4(_07813_),
    .ZN(_08104_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16233_ (.A1(_07981_),
    .A2(_08035_),
    .B1(_08009_),
    .B2(_07807_),
    .ZN(_08105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16234_ (.A1(_08104_),
    .A2(_08105_),
    .ZN(_08106_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16235_ (.A1(_08103_),
    .A2(_08106_),
    .Z(_08107_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16236_ (.A1(_08100_),
    .A2(_08107_),
    .ZN(_08108_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16237_ (.A1(_08099_),
    .A2(_08108_),
    .ZN(_08109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16238_ (.A1(_08080_),
    .A2(_08089_),
    .ZN(_08110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16239_ (.A1(_08080_),
    .A2(_08089_),
    .ZN(_08111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16240_ (.A1(_08079_),
    .A2(_08110_),
    .B(_08111_),
    .ZN(_08112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16241_ (.A1(_08109_),
    .A2(_08112_),
    .Z(_08113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16242_ (.A1(_08098_),
    .A2(_08113_),
    .ZN(_08114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16243_ (.A1(_08098_),
    .A2(_08113_),
    .ZN(_08115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16244_ (.A1(_07748_),
    .A2(_08115_),
    .ZN(_08116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16245_ (.I(_07749_),
    .Z(_08117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _16246_ (.A1(\spi_dac_i.spi_dat_buff_1[8] ),
    .A2(_07855_),
    .B1(_08114_),
    .B2(_08116_),
    .C(_08117_),
    .ZN(_08118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16247_ (.I(_07715_),
    .Z(_08119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16248_ (.A1(\spi_dac_i.spi_dat_buff_1[9] ),
    .A2(_07945_),
    .B(_08119_),
    .ZN(_08120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16249_ (.A1(_08118_),
    .A2(_08120_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16250_ (.A1(_08109_),
    .A2(_08112_),
    .ZN(_08121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16251_ (.A1(_08098_),
    .A2(_08113_),
    .B(_08121_),
    .ZN(_08122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16252_ (.A1(_08099_),
    .A2(_08108_),
    .ZN(_08123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16253_ (.A1(_08100_),
    .A2(_08107_),
    .B(_08123_),
    .ZN(_08124_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16254_ (.A1(_08103_),
    .A2(_08106_),
    .Z(_08125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16255_ (.A1(_08104_),
    .A2(_08125_),
    .ZN(_08126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16256_ (.A1(_08124_),
    .A2(_08126_),
    .Z(_08127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16257_ (.A1(_08122_),
    .A2(_08127_),
    .B(_07762_),
    .ZN(_08128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16258_ (.A1(_08122_),
    .A2(_08127_),
    .B(_08128_),
    .ZN(_08129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _16259_ (.A1(\spi_dac_i.spi_dat_buff_1[9] ),
    .A2(_07855_),
    .B(_08117_),
    .C(_08129_),
    .ZN(_08130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16260_ (.A1(\spi_dac_i.spi_dat_buff_1[10] ),
    .A2(_07891_),
    .B(_08119_),
    .ZN(_08131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16261_ (.A1(_08130_),
    .A2(_08131_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16262_ (.A1(_08104_),
    .A2(_08125_),
    .B(_08124_),
    .ZN(_08132_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16263_ (.A1(\spi_dac_i.spi_dat_buff_1[10] ),
    .A2(_07743_),
    .B1(_08132_),
    .B2(_08128_),
    .ZN(_08133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16264_ (.I(_07687_),
    .Z(_08134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16265_ (.A1(\spi_dac_i.spi_dat_buff_1[11] ),
    .A2(_07891_),
    .B(_08134_),
    .ZN(_08135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16266_ (.A1(_07945_),
    .A2(_08133_),
    .B(_08135_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16267_ (.A1(\filters.sample_buff[3] ),
    .A2(_07743_),
    .B1(_07750_),
    .B2(\spi_dac_i.spi_dat_buff_0[0] ),
    .ZN(_08136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16268_ (.A1(_07944_),
    .A2(_08136_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16269_ (.I(_07762_),
    .Z(_08137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16270_ (.A1(_07741_),
    .A2(_07738_),
    .ZN(_08138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16271_ (.I(_08138_),
    .Z(_08139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _16272_ (.A1(\filters.sample_buff[4] ),
    .A2(_08137_),
    .B1(_08139_),
    .B2(\spi_dac_i.spi_dat_buff_0[0] ),
    .C1(\spi_dac_i.spi_dat_buff_0[1] ),
    .C2(_07750_),
    .ZN(_08140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16273_ (.A1(_07944_),
    .A2(_08140_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16274_ (.I(_07749_),
    .Z(_08141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16275_ (.A1(\filters.sample_buff[5] ),
    .A2(_08137_),
    .B1(_08139_),
    .B2(\spi_dac_i.spi_dat_buff_0[1] ),
    .C1(\spi_dac_i.spi_dat_buff_0[2] ),
    .C2(_08141_),
    .ZN(_08142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16276_ (.A1(_07944_),
    .A2(_08142_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16277_ (.I(_07616_),
    .Z(_08143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16278_ (.I(_08138_),
    .Z(_08144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16279_ (.A1(\filters.sample_buff[6] ),
    .A2(_08137_),
    .B1(_08144_),
    .B2(\spi_dac_i.spi_dat_buff_0[2] ),
    .C1(\spi_dac_i.spi_dat_buff_0[3] ),
    .C2(_08141_),
    .ZN(_08145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16280_ (.A1(_08143_),
    .A2(_08145_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16281_ (.A1(\filters.sample_buff[7] ),
    .A2(_08137_),
    .B1(_08144_),
    .B2(\spi_dac_i.spi_dat_buff_0[3] ),
    .C1(\spi_dac_i.spi_dat_buff_0[4] ),
    .C2(_08141_),
    .ZN(_08146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16282_ (.A1(_08143_),
    .A2(_08146_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16283_ (.I(_07762_),
    .Z(_08147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16284_ (.A1(\filters.sample_buff[8] ),
    .A2(_08147_),
    .B1(_08144_),
    .B2(\spi_dac_i.spi_dat_buff_0[4] ),
    .C1(\spi_dac_i.spi_dat_buff_0[5] ),
    .C2(_08141_),
    .ZN(_08148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16285_ (.A1(_08143_),
    .A2(_08148_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16286_ (.I(_07749_),
    .Z(_08149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16287_ (.A1(\filters.sample_buff[9] ),
    .A2(_08147_),
    .B1(_08144_),
    .B2(\spi_dac_i.spi_dat_buff_0[5] ),
    .C1(\spi_dac_i.spi_dat_buff_0[6] ),
    .C2(_08149_),
    .ZN(_08150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16288_ (.A1(_08143_),
    .A2(_08150_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16289_ (.I(_07616_),
    .Z(_08151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16290_ (.I(_08138_),
    .Z(_08152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16291_ (.A1(\filters.sample_buff[10] ),
    .A2(_08147_),
    .B1(_08152_),
    .B2(\spi_dac_i.spi_dat_buff_0[6] ),
    .C1(\spi_dac_i.spi_dat_buff_0[7] ),
    .C2(_08149_),
    .ZN(_08153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16292_ (.A1(_08151_),
    .A2(_08153_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16293_ (.A1(\filters.sample_buff[11] ),
    .A2(_08147_),
    .B1(_08152_),
    .B2(\spi_dac_i.spi_dat_buff_0[7] ),
    .C1(\spi_dac_i.spi_dat_buff_0[8] ),
    .C2(_08149_),
    .ZN(_08154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16294_ (.A1(_08151_),
    .A2(_08154_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16295_ (.A1(\filters.sample_buff[12] ),
    .A2(_07763_),
    .B1(_08152_),
    .B2(\spi_dac_i.spi_dat_buff_0[8] ),
    .C1(\spi_dac_i.spi_dat_buff_0[9] ),
    .C2(_08149_),
    .ZN(_08155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16296_ (.A1(_08151_),
    .A2(_08155_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _16297_ (.A1(\filters.sample_buff[13] ),
    .A2(_07763_),
    .B1(_08152_),
    .B2(\spi_dac_i.spi_dat_buff_0[9] ),
    .C1(\spi_dac_i.spi_dat_buff_0[10] ),
    .C2(_08117_),
    .ZN(_08156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16298_ (.A1(_08151_),
    .A2(_08156_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16299_ (.I(_01943_),
    .Z(_08157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16300_ (.I(_08157_),
    .Z(_08158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _16301_ (.A1(\filters.sample_buff[14] ),
    .A2(_07763_),
    .B1(_08138_),
    .B2(\spi_dac_i.spi_dat_buff_0[10] ),
    .C1(\spi_dac_i.spi_dat_buff_0[11] ),
    .C2(_08117_),
    .ZN(_08159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16302_ (.A1(_08158_),
    .A2(_08159_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16303_ (.A1(net19),
    .A2(_07740_),
    .ZN(_08160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16304_ (.A1(\spi_dac_i.spi_dat_buff_1[11] ),
    .A2(_08139_),
    .ZN(_08161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16305_ (.A1(_08160_),
    .A2(_08161_),
    .B(_07745_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16306_ (.A1(net18),
    .A2(_07740_),
    .ZN(_08162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16307_ (.A1(\spi_dac_i.spi_dat_buff_0[11] ),
    .A2(_08139_),
    .ZN(_08163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16308_ (.A1(_08162_),
    .A2(_08163_),
    .B(_07745_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16309_ (.A1(_03510_),
    .A2(_07859_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16310_ (.A1(_03765_),
    .A2(_03769_),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16311_ (.A1(_02356_),
    .A2(_03770_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16312_ (.I(\channels.env_counter[3][0] ),
    .Z(_08164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16313_ (.I(_08164_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16314_ (.I(\channels.env_counter[3][1] ),
    .Z(_08165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16315_ (.I(_08165_),
    .Z(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16316_ (.I(\channels.env_counter[3][2] ),
    .Z(_08166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16317_ (.I(_08166_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16318_ (.I(\channels.env_counter[3][3] ),
    .Z(_08167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16319_ (.I(_08167_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16320_ (.I(\channels.env_counter[3][4] ),
    .Z(_08168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16321_ (.I(_08168_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16322_ (.I(\channels.env_counter[3][5] ),
    .Z(_08169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16323_ (.I(_08169_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16324_ (.I(\channels.env_counter[3][6] ),
    .Z(_08170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16325_ (.I(_08170_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16326_ (.I(\channels.env_counter[3][7] ),
    .Z(_08171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16327_ (.I(_08171_),
    .Z(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16328_ (.I(\channels.env_counter[3][8] ),
    .Z(_08172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16329_ (.I(_08172_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16330_ (.I(\channels.env_counter[3][9] ),
    .Z(_08173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16331_ (.I(_08173_),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16332_ (.I(\channels.env_counter[3][10] ),
    .Z(_08174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16333_ (.I(_08174_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16334_ (.I(\channels.env_counter[3][11] ),
    .Z(_08175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16335_ (.I(_08175_),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16336_ (.I(\channels.env_counter[3][12] ),
    .Z(_08176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16337_ (.I(_08176_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16338_ (.I(\channels.env_counter[3][13] ),
    .Z(_08177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16339_ (.I(_08177_),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16340_ (.I(\channels.env_counter[3][14] ),
    .Z(_08178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16341_ (.I(_08178_),
    .Z(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16342_ (.A1(_02365_),
    .A2(_03966_),
    .ZN(_08179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16343_ (.I(_08179_),
    .Z(_08180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16344_ (.A1(_02365_),
    .A2(_03965_),
    .B(_03650_),
    .ZN(_08181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16345_ (.I(_08181_),
    .Z(_08182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16346_ (.A1(\channels.env_vol[1][0] ),
    .A2(_08182_),
    .ZN(_08183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16347_ (.A1(_03772_),
    .A2(_08180_),
    .B(_08183_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16348_ (.A1(\channels.env_vol[1][1] ),
    .A2(_08182_),
    .ZN(_08184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16349_ (.A1(_03976_),
    .A2(_08180_),
    .B(_08184_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16350_ (.A1(\channels.env_vol[1][2] ),
    .A2(_08182_),
    .ZN(_08185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16351_ (.A1(_03982_),
    .A2(_08180_),
    .B(_08185_),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16352_ (.A1(\channels.env_vol[1][3] ),
    .A2(_08182_),
    .ZN(_08186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16353_ (.A1(_03986_),
    .A2(_08180_),
    .B(_08186_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16354_ (.I(_08179_),
    .Z(_08187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16355_ (.I(_08181_),
    .Z(_08188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16356_ (.A1(\channels.env_vol[1][4] ),
    .A2(_08188_),
    .ZN(_08189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16357_ (.A1(_03992_),
    .A2(_08187_),
    .B(_08189_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16358_ (.A1(\channels.env_vol[1][5] ),
    .A2(_08188_),
    .ZN(_08190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16359_ (.A1(_04002_),
    .A2(_08187_),
    .B(_08190_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16360_ (.A1(\channels.env_vol[1][6] ),
    .A2(_08188_),
    .ZN(_08191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16361_ (.A1(_04006_),
    .A2(_08187_),
    .B(_08191_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16362_ (.A1(\channels.env_vol[1][7] ),
    .A2(_08188_),
    .ZN(_08192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16363_ (.A1(_04009_),
    .A2(_08187_),
    .B(_08192_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16364_ (.A1(_01228_),
    .A2(_01265_),
    .B1(_01268_),
    .B2(\channels.exp_counter[0][0] ),
    .ZN(_08193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16365_ (.I(_08193_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16366_ (.A1(_01235_),
    .A2(_01265_),
    .B1(_01268_),
    .B2(\channels.exp_counter[0][1] ),
    .ZN(_08194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16367_ (.I(_08194_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16368_ (.A1(_01238_),
    .A2(_01327_),
    .B1(_01268_),
    .B2(\channels.exp_counter[0][2] ),
    .ZN(_08195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16369_ (.I(_08195_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16370_ (.A1(_01245_),
    .A2(_01327_),
    .B1(_01344_),
    .B2(\channels.exp_counter[0][3] ),
    .ZN(_08196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16371_ (.I(_08196_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16372_ (.A1(_01248_),
    .A2(_01327_),
    .B1(_01344_),
    .B2(\channels.exp_counter[0][4] ),
    .ZN(_08197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16373_ (.I(_08197_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16374_ (.A1(_02358_),
    .A2(_03966_),
    .ZN(_08198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16375_ (.I(_08198_),
    .Z(_08199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16376_ (.A1(_02358_),
    .A2(_03965_),
    .B(_01826_),
    .ZN(_08200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16377_ (.I(_08200_),
    .Z(_08201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16378_ (.A1(\channels.ch3_env[0] ),
    .A2(_08201_),
    .ZN(_08202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16379_ (.A1(_03772_),
    .A2(_08199_),
    .B(_08202_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16380_ (.A1(\channels.ch3_env[1] ),
    .A2(_08201_),
    .ZN(_08203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16381_ (.A1(_03976_),
    .A2(_08199_),
    .B(_08203_),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16382_ (.A1(\channels.ch3_env[2] ),
    .A2(_08201_),
    .ZN(_08204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16383_ (.A1(_03982_),
    .A2(_08199_),
    .B(_08204_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16384_ (.A1(\channels.ch3_env[3] ),
    .A2(_08201_),
    .ZN(_08205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16385_ (.A1(_03986_),
    .A2(_08199_),
    .B(_08205_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16386_ (.I(_08198_),
    .Z(_08206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16387_ (.I(_08200_),
    .Z(_08207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16388_ (.A1(\channels.ch3_env[4] ),
    .A2(_08207_),
    .ZN(_08208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16389_ (.A1(_03992_),
    .A2(_08206_),
    .B(_08208_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16390_ (.A1(\channels.ch3_env[5] ),
    .A2(_08207_),
    .ZN(_08209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16391_ (.A1(_04002_),
    .A2(_08206_),
    .B(_08209_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16392_ (.A1(\channels.ch3_env[6] ),
    .A2(_08207_),
    .ZN(_08210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16393_ (.A1(_04006_),
    .A2(_08206_),
    .B(_08210_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16394_ (.A1(\channels.ch3_env[7] ),
    .A2(_08207_),
    .ZN(_08211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16395_ (.A1(_04009_),
    .A2(_08206_),
    .B(_08211_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16396_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ),
    .A2(_02351_),
    .Z(_08212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16397_ (.I(_08212_),
    .Z(_08213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16398_ (.I(_08213_),
    .Z(_08214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16399_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ),
    .A2(_08213_),
    .ZN(_08215_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _16400_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.restart_noise ),
    .A2(_01040_),
    .Z(_08216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16401_ (.I(_08216_),
    .Z(_08217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _16402_ (.A1(_07830_),
    .A2(_08214_),
    .B(_08215_),
    .C(_08217_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16403_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ),
    .A2(_08214_),
    .ZN(_08218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16404_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ),
    .A2(_02351_),
    .ZN(_08219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16405_ (.I(_08219_),
    .Z(_08220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16406_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ),
    .A2(_08220_),
    .ZN(_08221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16407_ (.I(_08217_),
    .Z(_08222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16408_ (.A1(_08218_),
    .A2(_08221_),
    .B(_08222_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16409_ (.I(_08213_),
    .Z(_08223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16410_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ),
    .A2(_08223_),
    .ZN(_08224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16411_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ),
    .A2(_08220_),
    .ZN(_08225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16412_ (.A1(_08224_),
    .A2(_08225_),
    .B(_08222_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16413_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ),
    .A2(_08223_),
    .ZN(_08226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16414_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ),
    .A2(_08220_),
    .ZN(_08227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16415_ (.A1(_08226_),
    .A2(_08227_),
    .B(_08222_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16416_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ),
    .A2(_08223_),
    .ZN(_08228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16417_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ),
    .A2(_08220_),
    .ZN(_08229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16418_ (.A1(_08228_),
    .A2(_08229_),
    .B(_08222_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16419_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ),
    .A2(_08223_),
    .ZN(_08230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16420_ (.I(_08219_),
    .Z(_08231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16421_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ),
    .A2(_08231_),
    .ZN(_08232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16422_ (.I(_08216_),
    .Z(_08233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16423_ (.A1(_08230_),
    .A2(_08232_),
    .B(_08233_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16424_ (.I(_08213_),
    .Z(_08234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16425_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ),
    .A2(_08234_),
    .ZN(_08235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16426_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ),
    .A2(_08231_),
    .ZN(_08236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16427_ (.A1(_08235_),
    .A2(_08236_),
    .B(_08233_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16428_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ),
    .A2(_08234_),
    .ZN(_08237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16429_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ),
    .A2(_08231_),
    .ZN(_08238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16430_ (.A1(_08237_),
    .A2(_08238_),
    .B(_08233_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16431_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ),
    .A2(_08234_),
    .ZN(_08239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16432_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ),
    .A2(_08231_),
    .ZN(_08240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16433_ (.A1(_08239_),
    .A2(_08240_),
    .B(_08233_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16434_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ),
    .A2(_08234_),
    .ZN(_08241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16435_ (.I(_08219_),
    .Z(_08242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16436_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ),
    .A2(_08242_),
    .ZN(_08243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16437_ (.I(_08216_),
    .Z(_08244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16438_ (.A1(_08241_),
    .A2(_08243_),
    .B(_08244_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16439_ (.I(_08212_),
    .Z(_08245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16440_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ),
    .A2(_08245_),
    .ZN(_08246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16441_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ),
    .A2(_08242_),
    .ZN(_08247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16442_ (.A1(_08246_),
    .A2(_08247_),
    .B(_08244_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16443_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ),
    .A2(_08245_),
    .ZN(_08248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16444_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ),
    .A2(_08242_),
    .ZN(_08249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16445_ (.A1(_08248_),
    .A2(_08249_),
    .B(_08244_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16446_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ),
    .A2(_08245_),
    .ZN(_08250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16447_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ),
    .A2(_08242_),
    .ZN(_08251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16448_ (.A1(_08250_),
    .A2(_08251_),
    .B(_08244_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16449_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ),
    .A2(_08245_),
    .ZN(_08252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16450_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ),
    .A2(_08219_),
    .ZN(_08253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16451_ (.A1(_08252_),
    .A2(_08253_),
    .B(_08217_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16452_ (.A1(\tt_um_rejunity_sn76489.control_noise[0][2] ),
    .A2(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ),
    .ZN(_08254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16453_ (.A1(_07839_),
    .A2(_08254_),
    .Z(_08255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16454_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ),
    .A2(_08214_),
    .B(_08217_),
    .ZN(_08256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16455_ (.A1(_08214_),
    .A2(_08255_),
    .B(_08256_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16456_ (.A1(\tt_um_rejunity_sn76489.clk_counter[4] ),
    .A2(\tt_um_rejunity_sn76489.clk_counter[3] ),
    .ZN(_08257_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _16457_ (.A1(\tt_um_rejunity_sn76489.clk_counter[2] ),
    .A2(\tt_um_rejunity_sn76489.clk_counter[1] ),
    .A3(\tt_um_rejunity_sn76489.clk_counter[0] ),
    .ZN(_08258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16458_ (.A1(_08257_),
    .A2(_08258_),
    .ZN(_08259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16459_ (.I(_08259_),
    .Z(_08260_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16460_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[0] ),
    .A2(_08260_),
    .Z(_08261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16461_ (.A1(_08158_),
    .A2(_08261_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16462_ (.A1(_08257_),
    .A2(_08258_),
    .Z(_08262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16463_ (.I(_08262_),
    .Z(_08263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16464_ (.I(_08263_),
    .Z(_08264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16465_ (.I(_08264_),
    .Z(_08265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16466_ (.I(_08265_),
    .Z(_08266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16467_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[0] ),
    .A2(_08266_),
    .B(\tt_um_rejunity_sn76489.noise[0].gen.counter[1] ),
    .ZN(_08267_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16468_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[1] ),
    .A2(\tt_um_rejunity_sn76489.noise[0].gen.counter[0] ),
    .A3(_08262_),
    .Z(_08268_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16469_ (.A1(_04129_),
    .A2(_08267_),
    .A3(_08268_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16470_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[2] ),
    .A2(_08268_),
    .Z(_08269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16471_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[2] ),
    .A2(_08268_),
    .B(_08119_),
    .ZN(_08270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16472_ (.A1(_08269_),
    .A2(_08270_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16473_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[3] ),
    .A2(_08269_),
    .Z(_08271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16474_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[3] ),
    .A2(_08269_),
    .B(_08119_),
    .ZN(_08272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16475_ (.A1(_08271_),
    .A2(_08272_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16476_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ),
    .A2(_08271_),
    .Z(_08273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16477_ (.I(_07715_),
    .Z(_08274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16478_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ),
    .A2(_08271_),
    .B(_08274_),
    .ZN(_08275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16479_ (.A1(_08273_),
    .A2(_08275_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16480_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ),
    .A2(_08273_),
    .B(_08134_),
    .ZN(_08276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16481_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ),
    .A2(_08273_),
    .B(_08276_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16482_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ),
    .A2(_08273_),
    .ZN(_08277_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16483_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.counter[6] ),
    .A2(_08277_),
    .Z(_08278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16484_ (.A1(_08158_),
    .A2(_08278_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16485_ (.A1(_08158_),
    .A2(_07945_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16486_ (.I(_08263_),
    .Z(_08279_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16487_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ),
    .A2(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ),
    .A3(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ),
    .A4(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ),
    .Z(_08280_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16488_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ),
    .A2(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ),
    .A3(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ),
    .A4(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ),
    .Z(_08281_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _16489_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[9] ),
    .A2(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ),
    .A3(_08280_),
    .A4(_08281_),
    .ZN(_08282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16490_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][0] ),
    .A2(_08282_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ),
    .ZN(_08283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16491_ (.A1(_08279_),
    .A2(_08283_),
    .ZN(_08284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16492_ (.I(_08259_),
    .Z(_08285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16493_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ),
    .A2(_08285_),
    .ZN(_08286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16494_ (.I(_07566_),
    .Z(_08287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16495_ (.A1(_08284_),
    .A2(_08286_),
    .B(_08287_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16496_ (.I(_08157_),
    .Z(_08288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16497_ (.I(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ),
    .ZN(_08289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16498_ (.I(_08263_),
    .Z(_08290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16499_ (.I(_08282_),
    .Z(_08291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16500_ (.I(_08291_),
    .Z(_08292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16501_ (.I(_08292_),
    .Z(_08293_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16502_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ),
    .A2(_08290_),
    .A3(_08293_),
    .ZN(_08294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16503_ (.A1(_08289_),
    .A2(_08294_),
    .ZN(_08295_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16504_ (.A1(_08284_),
    .A2(_08295_),
    .Z(_08296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16505_ (.A1(_08288_),
    .A2(_08296_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16506_ (.I(_08259_),
    .Z(_08297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16507_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][2] ),
    .A2(_08291_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ),
    .ZN(_08298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16508_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ),
    .A2(_08291_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ),
    .ZN(_08299_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16509_ (.A1(_08283_),
    .A2(_08298_),
    .A3(_08299_),
    .Z(_08300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16510_ (.A1(_08283_),
    .A2(_08299_),
    .B(_08298_),
    .ZN(_08301_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16511_ (.A1(_08297_),
    .A2(_08300_),
    .A3(_08301_),
    .ZN(_08302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16512_ (.I(_08263_),
    .Z(_08303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16513_ (.I(_08303_),
    .Z(_08304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16514_ (.I(_08304_),
    .Z(_08305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16515_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ),
    .A2(_08305_),
    .B(_08274_),
    .ZN(_08306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16516_ (.A1(_08302_),
    .A2(_08306_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16517_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][3] ),
    .A2(_08291_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ),
    .ZN(_08307_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16518_ (.A1(_08300_),
    .A2(_08307_),
    .Z(_08308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16519_ (.A1(_08300_),
    .A2(_08307_),
    .B(_08266_),
    .ZN(_08309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16520_ (.A1(_08308_),
    .A2(_08309_),
    .ZN(_08310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16521_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ),
    .A2(_08305_),
    .B(_08274_),
    .ZN(_08311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16522_ (.A1(_08310_),
    .A2(_08311_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16523_ (.I(_08265_),
    .Z(_08312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16524_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][4] ),
    .A2(_08292_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ),
    .ZN(_08313_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16525_ (.A1(_08308_),
    .A2(_08313_),
    .Z(_08314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16526_ (.I(_08279_),
    .Z(_08315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16527_ (.A1(_08308_),
    .A2(_08313_),
    .B(_08315_),
    .ZN(_08316_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16528_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ),
    .A2(_08312_),
    .B1(_08314_),
    .B2(_08316_),
    .ZN(_08317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16529_ (.A1(_08288_),
    .A2(_08317_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16530_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][5] ),
    .A2(_08292_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ),
    .ZN(_08318_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16531_ (.A1(_08314_),
    .A2(_08318_),
    .Z(_08319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16532_ (.A1(_08314_),
    .A2(_08318_),
    .B(_08315_),
    .ZN(_08320_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16533_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ),
    .A2(_08312_),
    .B1(_08319_),
    .B2(_08320_),
    .ZN(_08321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16534_ (.A1(_08288_),
    .A2(_08321_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16535_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][6] ),
    .A2(_08292_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ),
    .ZN(_08322_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16536_ (.A1(_08319_),
    .A2(_08322_),
    .Z(_08323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16537_ (.I(_08279_),
    .Z(_08324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16538_ (.A1(_08319_),
    .A2(_08322_),
    .B(_08324_),
    .ZN(_08325_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16539_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ),
    .A2(_08312_),
    .B1(_08323_),
    .B2(_08325_),
    .ZN(_08326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16540_ (.A1(_08288_),
    .A2(_08326_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16541_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][7] ),
    .A2(_08293_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ),
    .ZN(_08327_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16542_ (.A1(_08323_),
    .A2(_08327_),
    .Z(_08328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16543_ (.A1(_08323_),
    .A2(_08327_),
    .ZN(_08329_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16544_ (.A1(_08297_),
    .A2(_08328_),
    .A3(_08329_),
    .ZN(_08330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16545_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ),
    .A2(_08305_),
    .B(_08274_),
    .ZN(_08331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16546_ (.A1(_08330_),
    .A2(_08331_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16547_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][8] ),
    .A2(_08293_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ),
    .ZN(_08332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16548_ (.A1(_08303_),
    .A2(_08328_),
    .A3(_08332_),
    .ZN(_08333_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16549_ (.A1(_08260_),
    .A2(_08328_),
    .A3(_08332_),
    .ZN(_08334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16550_ (.A1(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ),
    .A2(_08285_),
    .B(_08334_),
    .ZN(_08335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16551_ (.A1(_08333_),
    .A2(_08335_),
    .B(_08287_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16552_ (.I(_08157_),
    .Z(_08336_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16553_ (.A1(_08264_),
    .A2(_08293_),
    .Z(_08337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16554_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][9] ),
    .A2(_08337_),
    .B(\tt_um_rejunity_sn76489.tone[2].gen.counter[9] ),
    .ZN(_08338_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16555_ (.A1(_08333_),
    .A2(_08338_),
    .ZN(_08339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16556_ (.A1(_08336_),
    .A2(_08339_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16557_ (.A1(_02349_),
    .A2(_08337_),
    .B(_08134_),
    .ZN(_08340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16558_ (.A1(_02349_),
    .A2(_08337_),
    .B(_08340_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16559_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ),
    .A2(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ),
    .A3(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ),
    .A4(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ),
    .Z(_08341_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16560_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ),
    .A2(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ),
    .A3(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ),
    .A4(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ),
    .Z(_08342_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _16561_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[9] ),
    .A2(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ),
    .A3(_08341_),
    .A4(_08342_),
    .ZN(_08343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16562_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][0] ),
    .A2(_08343_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ),
    .ZN(_08344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16563_ (.A1(_08279_),
    .A2(_08344_),
    .ZN(_08345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16564_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ),
    .A2(_08285_),
    .ZN(_08346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16565_ (.A1(_08345_),
    .A2(_08346_),
    .B(_08287_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16566_ (.I(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ),
    .ZN(_08347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16567_ (.I(_08343_),
    .Z(_08348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16568_ (.I(_08348_),
    .Z(_08349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16569_ (.I(_08349_),
    .Z(_08350_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16570_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ),
    .A2(_08290_),
    .A3(_08350_),
    .ZN(_08351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16571_ (.A1(_08347_),
    .A2(_08351_),
    .ZN(_08352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16572_ (.A1(_08345_),
    .A2(_08352_),
    .Z(_08353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16573_ (.A1(_08336_),
    .A2(_08353_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16574_ (.I(_08259_),
    .Z(_08354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16575_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][2] ),
    .A2(_08348_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ),
    .ZN(_08355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16576_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ),
    .A2(_08348_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ),
    .ZN(_08356_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16577_ (.A1(_08344_),
    .A2(_08355_),
    .A3(_08356_),
    .Z(_08357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16578_ (.A1(_08344_),
    .A2(_08356_),
    .B(_08355_),
    .ZN(_08358_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16579_ (.A1(_08354_),
    .A2(_08357_),
    .A3(_08358_),
    .ZN(_08359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16580_ (.I(_07715_),
    .Z(_08360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16581_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ),
    .A2(_08305_),
    .B(_08360_),
    .ZN(_08361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16582_ (.A1(_08359_),
    .A2(_08361_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16583_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][3] ),
    .A2(_08348_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ),
    .ZN(_08362_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16584_ (.A1(_08357_),
    .A2(_08362_),
    .Z(_08363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16585_ (.A1(_08357_),
    .A2(_08362_),
    .B(_08315_),
    .ZN(_08364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16586_ (.A1(_08363_),
    .A2(_08364_),
    .ZN(_08365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16587_ (.I(_08265_),
    .Z(_08366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16588_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ),
    .A2(_08366_),
    .B(_08360_),
    .ZN(_08367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16589_ (.A1(_08365_),
    .A2(_08367_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16590_ (.I(_08265_),
    .Z(_08368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16591_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][4] ),
    .A2(_08349_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ),
    .ZN(_08369_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16592_ (.A1(_08363_),
    .A2(_08369_),
    .Z(_08370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16593_ (.A1(_08363_),
    .A2(_08369_),
    .B(_08324_),
    .ZN(_08371_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16594_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ),
    .A2(_08368_),
    .B1(_08370_),
    .B2(_08371_),
    .ZN(_08372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16595_ (.A1(_08336_),
    .A2(_08372_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16596_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][5] ),
    .A2(_08349_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ),
    .ZN(_08373_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16597_ (.A1(_08370_),
    .A2(_08373_),
    .Z(_08374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16598_ (.A1(_08370_),
    .A2(_08373_),
    .B(_08324_),
    .ZN(_08375_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16599_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ),
    .A2(_08368_),
    .B1(_08374_),
    .B2(_08375_),
    .ZN(_08376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16600_ (.A1(_08336_),
    .A2(_08376_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16601_ (.I(_08157_),
    .Z(_08377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16602_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][6] ),
    .A2(_08349_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ),
    .ZN(_08378_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16603_ (.A1(_08374_),
    .A2(_08378_),
    .Z(_08379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16604_ (.A1(_08374_),
    .A2(_08378_),
    .B(_08324_),
    .ZN(_08380_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16605_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ),
    .A2(_08368_),
    .B1(_08379_),
    .B2(_08380_),
    .ZN(_08381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16606_ (.A1(_08377_),
    .A2(_08381_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16607_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][7] ),
    .A2(_08350_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ),
    .ZN(_08382_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16608_ (.A1(_08379_),
    .A2(_08382_),
    .Z(_08383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16609_ (.A1(_08379_),
    .A2(_08382_),
    .ZN(_08384_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16610_ (.A1(_08354_),
    .A2(_08383_),
    .A3(_08384_),
    .ZN(_08385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16611_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ),
    .A2(_08366_),
    .B(_08360_),
    .ZN(_08386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16612_ (.A1(_08385_),
    .A2(_08386_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16613_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][8] ),
    .A2(_08350_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ),
    .ZN(_08387_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16614_ (.A1(_08303_),
    .A2(_08383_),
    .A3(_08387_),
    .ZN(_08388_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16615_ (.A1(_08260_),
    .A2(_08383_),
    .A3(_08387_),
    .ZN(_08389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16616_ (.A1(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ),
    .A2(_08297_),
    .B(_08389_),
    .ZN(_08390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16617_ (.A1(_08388_),
    .A2(_08390_),
    .B(_08287_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16618_ (.A1(_08264_),
    .A2(_08350_),
    .Z(_08391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16619_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][9] ),
    .A2(_08391_),
    .B(\tt_um_rejunity_sn76489.tone[1].gen.counter[9] ),
    .ZN(_08392_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16620_ (.A1(_08388_),
    .A2(_08392_),
    .ZN(_08393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16621_ (.A1(_08377_),
    .A2(_08393_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16622_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.in ),
    .A2(_08391_),
    .B(_08134_),
    .ZN(_08394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16623_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.in ),
    .A2(_08391_),
    .B(_08394_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _16624_ (.A1(_01329_),
    .A2(_01597_),
    .Z(_08395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16625_ (.I(_08395_),
    .Z(_08396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16626_ (.I(_08396_),
    .Z(_08397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16627_ (.A1(_01600_),
    .A2(_08395_),
    .ZN(_08398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16628_ (.I(_08398_),
    .Z(_08399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16629_ (.I(_08399_),
    .Z(_08400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16630_ (.A1(_01590_),
    .A2(_08397_),
    .B1(_08400_),
    .B2(_01606_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16631_ (.A1(_01609_),
    .A2(_08397_),
    .B1(_08400_),
    .B2(_01612_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16632_ (.A1(_01619_),
    .A2(_08397_),
    .B1(_08400_),
    .B2(_01623_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16633_ (.A1(_01626_),
    .A2(_08397_),
    .B1(_08400_),
    .B2(_01628_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16634_ (.I(_08395_),
    .Z(_08401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16635_ (.I(_08401_),
    .Z(_08402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16636_ (.I(_08398_),
    .Z(_08403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16637_ (.I(_08403_),
    .Z(_08404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16638_ (.A1(_01631_),
    .A2(_08402_),
    .B1(_08404_),
    .B2(_01633_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16639_ (.A1(_01636_),
    .A2(_08402_),
    .B1(_08404_),
    .B2(_01640_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16640_ (.A1(_01643_),
    .A2(_08402_),
    .B1(_08404_),
    .B2(_01646_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16641_ (.A1(_01649_),
    .A2(_08402_),
    .B1(_08404_),
    .B2(_01651_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16642_ (.I(_08401_),
    .Z(_08405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16643_ (.I(_08403_),
    .Z(_08406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16644_ (.A1(_01656_),
    .A2(_08405_),
    .B1(_08406_),
    .B2(_01658_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16645_ (.A1(_01661_),
    .A2(_08405_),
    .B1(_08406_),
    .B2(_01664_),
    .ZN(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16646_ (.A1(_01668_),
    .A2(_08405_),
    .B1(_08406_),
    .B2(_01671_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16647_ (.A1(_01674_),
    .A2(_08405_),
    .B1(_08406_),
    .B2(_01676_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16648_ (.I(_08401_),
    .Z(_08407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16649_ (.I(_08403_),
    .Z(_08408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16650_ (.A1(_01679_),
    .A2(_08407_),
    .B1(_08408_),
    .B2(_01681_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16651_ (.A1(_01684_),
    .A2(_08407_),
    .B1(_08408_),
    .B2(_01687_),
    .ZN(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16652_ (.A1(_01692_),
    .A2(_08407_),
    .B1(_08408_),
    .B2(_01695_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16653_ (.A1(_01700_),
    .A2(_08407_),
    .B1(_08408_),
    .B2(_01702_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16654_ (.I(_08401_),
    .Z(_08409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16655_ (.I(_08403_),
    .Z(_08410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16656_ (.A1(_01705_),
    .A2(_08409_),
    .B1(_08410_),
    .B2(_01706_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16657_ (.A1(_01709_),
    .A2(_08409_),
    .B1(_08410_),
    .B2(_01583_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16658_ (.A1(_01587_),
    .A2(_08409_),
    .B1(_08410_),
    .B2(_01713_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16659_ (.A1(_01716_),
    .A2(_08409_),
    .B1(_08410_),
    .B2(_01718_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16660_ (.A1(_01721_),
    .A2(_08396_),
    .B1(_08399_),
    .B2(_01723_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16661_ (.A1(_01726_),
    .A2(_08396_),
    .B1(_08399_),
    .B2(_01728_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16662_ (.I(\channels.lfsr[0][22] ),
    .ZN(_08411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _16663_ (.A1(_01731_),
    .A2(_08396_),
    .B1(_08399_),
    .B2(_08411_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16664_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ),
    .A2(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ),
    .A3(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ),
    .A4(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ),
    .Z(_08412_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16665_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ),
    .A2(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ),
    .A3(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ),
    .A4(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ),
    .Z(_08413_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _16666_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[9] ),
    .A2(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ),
    .A3(_08412_),
    .A4(_08413_),
    .ZN(_08414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16667_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][0] ),
    .A2(_08414_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ),
    .ZN(_08415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16668_ (.A1(_08290_),
    .A2(_08415_),
    .ZN(_08416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16669_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ),
    .A2(_08285_),
    .ZN(_08417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16670_ (.I(_07566_),
    .Z(_08418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16671_ (.A1(_08416_),
    .A2(_08417_),
    .B(_08418_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16672_ (.I(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ),
    .ZN(_08419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16673_ (.I(_08414_),
    .Z(_08420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16674_ (.I(_08420_),
    .Z(_08421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16675_ (.I(_08421_),
    .Z(_08422_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16676_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][1] ),
    .A2(_08290_),
    .A3(_08422_),
    .ZN(_08423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16677_ (.A1(_08419_),
    .A2(_08423_),
    .ZN(_08424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16678_ (.A1(_08416_),
    .A2(_08424_),
    .Z(_08425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16679_ (.A1(_08377_),
    .A2(_08425_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16680_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][2] ),
    .A2(_08420_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ),
    .ZN(_08426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16681_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][1] ),
    .A2(_08420_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ),
    .ZN(_08427_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16682_ (.A1(_08415_),
    .A2(_08426_),
    .A3(_08427_),
    .Z(_08428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16683_ (.A1(_08415_),
    .A2(_08427_),
    .B(_08426_),
    .ZN(_08429_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16684_ (.A1(_08354_),
    .A2(_08428_),
    .A3(_08429_),
    .ZN(_08430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16685_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ),
    .A2(_08366_),
    .B(_08360_),
    .ZN(_08431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16686_ (.A1(_08430_),
    .A2(_08431_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16687_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][3] ),
    .A2(_08420_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ),
    .ZN(_08432_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16688_ (.A1(_08428_),
    .A2(_08432_),
    .Z(_08433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16689_ (.A1(_08428_),
    .A2(_08432_),
    .B(_08315_),
    .ZN(_08434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16690_ (.A1(_08433_),
    .A2(_08434_),
    .ZN(_08435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16691_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ),
    .A2(_08366_),
    .B(_01763_),
    .ZN(_08436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16692_ (.A1(_08435_),
    .A2(_08436_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16693_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][4] ),
    .A2(_08421_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ),
    .ZN(_08437_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16694_ (.A1(_08433_),
    .A2(_08437_),
    .Z(_08438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16695_ (.A1(_08433_),
    .A2(_08437_),
    .B(_08304_),
    .ZN(_08439_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16696_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ),
    .A2(_08368_),
    .B1(_08438_),
    .B2(_08439_),
    .ZN(_08440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16697_ (.A1(_08377_),
    .A2(_08440_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16698_ (.I(_03651_),
    .Z(_08441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16699_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][5] ),
    .A2(_08421_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ),
    .ZN(_08442_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16700_ (.A1(_08438_),
    .A2(_08442_),
    .Z(_08443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16701_ (.A1(_08438_),
    .A2(_08442_),
    .B(_08304_),
    .ZN(_08444_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16702_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ),
    .A2(_08266_),
    .B1(_08443_),
    .B2(_08444_),
    .ZN(_08445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16703_ (.A1(_08441_),
    .A2(_08445_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16704_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][6] ),
    .A2(_08421_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ),
    .ZN(_08446_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16705_ (.A1(_08443_),
    .A2(_08446_),
    .Z(_08447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16706_ (.A1(_08443_),
    .A2(_08446_),
    .B(_08304_),
    .ZN(_08448_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _16707_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ),
    .A2(_08266_),
    .B1(_08447_),
    .B2(_08448_),
    .ZN(_08449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16708_ (.A1(_08441_),
    .A2(_08449_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16709_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][7] ),
    .A2(_08422_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ),
    .ZN(_08450_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16710_ (.A1(_08447_),
    .A2(_08450_),
    .Z(_08451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16711_ (.A1(_08447_),
    .A2(_08450_),
    .ZN(_08452_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16712_ (.A1(_08354_),
    .A2(_08451_),
    .A3(_08452_),
    .ZN(_08453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16713_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ),
    .A2(_08312_),
    .B(_01763_),
    .ZN(_08454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16714_ (.A1(_08453_),
    .A2(_08454_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16715_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][8] ),
    .A2(_08422_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ),
    .ZN(_08455_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16716_ (.A1(_08303_),
    .A2(_08451_),
    .A3(_08455_),
    .ZN(_08456_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16717_ (.A1(_08260_),
    .A2(_08451_),
    .A3(_08455_),
    .ZN(_08457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16718_ (.A1(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ),
    .A2(_08297_),
    .B(_08457_),
    .ZN(_08458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16719_ (.A1(_08456_),
    .A2(_08458_),
    .B(_08418_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16720_ (.A1(_08264_),
    .A2(_08422_),
    .Z(_08459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16721_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][9] ),
    .A2(_08459_),
    .B(\tt_um_rejunity_sn76489.tone[0].gen.counter[9] ),
    .ZN(_08460_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _16722_ (.A1(_08456_),
    .A2(_08460_),
    .ZN(_08461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16723_ (.A1(_08441_),
    .A2(_08461_),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16724_ (.I(_07687_),
    .Z(_08462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16725_ (.A1(_07819_),
    .A2(_08459_),
    .B(_08462_),
    .ZN(_08463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16726_ (.A1(_07819_),
    .A2(_08459_),
    .B(_08463_),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16727_ (.I(\tt_um_rejunity_sn76489.latch_control_reg[2] ),
    .Z(_08464_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _16728_ (.A1(\tt_um_rejunity_sn76489.latch_control_reg[1] ),
    .A2(net14),
    .A3(_03497_),
    .ZN(_08465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16729_ (.A1(\tt_um_rejunity_sn76489.latch_control_reg[0] ),
    .A2(_03499_),
    .ZN(_08466_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16730_ (.A1(_08464_),
    .A2(_08465_),
    .A3(_08466_),
    .Z(_08467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16731_ (.I(_08467_),
    .Z(_08468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16732_ (.I(_08468_),
    .Z(_08469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16733_ (.I(_08467_),
    .Z(_08470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16734_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][4] ),
    .A2(_08470_),
    .B(_08462_),
    .ZN(_08471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16735_ (.A1(_03735_),
    .A2(_08469_),
    .B(_08471_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16736_ (.I(_01765_),
    .Z(_08472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16737_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][5] ),
    .A2(_08470_),
    .B(_08462_),
    .ZN(_08473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16738_ (.A1(_08472_),
    .A2(_08469_),
    .B(_08473_),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16739_ (.I(_01775_),
    .Z(_08474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16740_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][6] ),
    .A2(_08468_),
    .B(_08462_),
    .ZN(_08475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16741_ (.A1(_08474_),
    .A2(_08469_),
    .B(_08475_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16742_ (.I(_07687_),
    .Z(_08476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16743_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][7] ),
    .A2(_08468_),
    .B(_08476_),
    .ZN(_08477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16744_ (.A1(_03707_),
    .A2(_08469_),
    .B(_08477_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16745_ (.A1(_08464_),
    .A2(_08465_),
    .A3(_08466_),
    .ZN(_08478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16746_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][8] ),
    .A2(_08478_),
    .ZN(_08479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16747_ (.A1(_03747_),
    .A2(_08470_),
    .ZN(_08480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16748_ (.A1(_08479_),
    .A2(_08480_),
    .B(_08418_),
    .ZN(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16749_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[2][9] ),
    .A2(_08468_),
    .B(_08476_),
    .ZN(_08481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16750_ (.A1(_01811_),
    .A2(_08470_),
    .B(_08481_),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16751_ (.I(\tt_um_rejunity_sn76489.latch_control_reg[1] ),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16752_ (.A1(_03496_),
    .A2(_04186_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _16753_ (.A1(\tt_um_rejunity_sn76489.latch_control_reg[2] ),
    .A2(\tt_um_rejunity_sn76489.latch_control_reg[0] ),
    .A3(_03499_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16754_ (.A1(_00860_),
    .A2(_00861_),
    .A3(_00862_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16755_ (.I(_00863_),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16756_ (.I(_00864_),
    .Z(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16757_ (.I(_00863_),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16758_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][4] ),
    .A2(_00866_),
    .B(_08476_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16759_ (.A1(_03735_),
    .A2(_00865_),
    .B(_00867_),
    .ZN(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16760_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][5] ),
    .A2(_00866_),
    .B(_08476_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16761_ (.A1(_08472_),
    .A2(_00865_),
    .B(_00868_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16762_ (.I(_03766_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16763_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][6] ),
    .A2(_00864_),
    .B(_00869_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16764_ (.A1(_08474_),
    .A2(_00865_),
    .B(_00870_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16765_ (.I(_02320_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16766_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][7] ),
    .A2(_00864_),
    .B(_00869_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16767_ (.A1(_00871_),
    .A2(_00865_),
    .B(_00872_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16768_ (.A1(_00860_),
    .A2(_00861_),
    .A3(_00862_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16769_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][8] ),
    .A2(_00873_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16770_ (.A1(_03747_),
    .A2(_00866_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16771_ (.A1(_00874_),
    .A2(_00875_),
    .B(_08418_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16772_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[1][9] ),
    .A2(_00864_),
    .B(_00869_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16773_ (.A1(_01811_),
    .A2(_00866_),
    .B(_00876_),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16774_ (.A1(_08465_),
    .A2(_00862_),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16775_ (.I(_00877_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16776_ (.I(_00878_),
    .Z(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16777_ (.I(_00877_),
    .Z(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16778_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][4] ),
    .A2(_00880_),
    .B(_00869_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16779_ (.A1(_03735_),
    .A2(_00879_),
    .B(_00881_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16780_ (.I(_03766_),
    .Z(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16781_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][5] ),
    .A2(_00880_),
    .B(_00882_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16782_ (.A1(_08472_),
    .A2(_00879_),
    .B(_00883_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16783_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][6] ),
    .A2(_00878_),
    .B(_00882_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16784_ (.A1(_08474_),
    .A2(_00879_),
    .B(_00884_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16785_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][7] ),
    .A2(_00878_),
    .B(_00882_),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16786_ (.A1(_00871_),
    .A2(_00879_),
    .B(_00885_),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16787_ (.A1(_08465_),
    .A2(_00862_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16788_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][8] ),
    .A2(_00886_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16789_ (.A1(_03747_),
    .A2(_00880_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16790_ (.A1(_00887_),
    .A2(_00888_),
    .B(_01828_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16791_ (.A1(\tt_um_rejunity_sn76489.control_tone_freq[0][9] ),
    .A2(_00878_),
    .B(_00882_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16792_ (.A1(_01811_),
    .A2(_00880_),
    .B(_00889_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16793_ (.I(_03500_),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16794_ (.I(\tt_um_rejunity_sn76489.latch_control_reg[2] ),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16795_ (.I(\tt_um_rejunity_sn76489.latch_control_reg[1] ),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16796_ (.A1(\tt_um_rejunity_sn76489.latch_control_reg[0] ),
    .A2(_01820_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16797_ (.A1(_01815_),
    .A2(_03496_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16798_ (.A1(_03493_),
    .A2(_03494_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _16799_ (.A1(_00891_),
    .A2(_00892_),
    .A3(_00893_),
    .B1(_00894_),
    .B2(_00895_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16800_ (.A1(_00890_),
    .A2(_00896_),
    .Z(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16801_ (.I(_00897_),
    .Z(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16802_ (.I(_00897_),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16803_ (.A1(_03505_),
    .A2(_00899_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16804_ (.I(_03767_),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16805_ (.A1(_07847_),
    .A2(_00898_),
    .B(_00900_),
    .C(_00901_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16806_ (.A1(net8),
    .A2(_00899_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16807_ (.A1(_07842_),
    .A2(_00898_),
    .B(_00902_),
    .C(_00901_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16808_ (.A1(net9),
    .A2(_00899_),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16809_ (.A1(_07838_),
    .A2(_00898_),
    .B(_00903_),
    .C(_00901_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16810_ (.A1(net10),
    .A2(_00899_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16811_ (.A1(_07930_),
    .A2(_00898_),
    .B(_00904_),
    .C(_00901_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16812_ (.I(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16813_ (.A1(_01042_),
    .A2(_03494_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _16814_ (.A1(_00891_),
    .A2(_00860_),
    .A3(_00893_),
    .B1(_00906_),
    .B2(_00894_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16815_ (.A1(_03500_),
    .A2(_00907_),
    .Z(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16816_ (.I(_00908_),
    .Z(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16817_ (.I(_00908_),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16818_ (.A1(_03505_),
    .A2(_00910_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16819_ (.I(_03767_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16820_ (.A1(_00905_),
    .A2(_00909_),
    .B(_00911_),
    .C(_00912_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16821_ (.I(_07862_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16822_ (.A1(net8),
    .A2(_00910_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16823_ (.A1(_00913_),
    .A2(_00909_),
    .B(_00914_),
    .C(_00912_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16824_ (.A1(net9),
    .A2(_00910_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16825_ (.A1(_07776_),
    .A2(_00909_),
    .B(_00915_),
    .C(_00912_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16826_ (.A1(net10),
    .A2(_00910_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16827_ (.A1(_07780_),
    .A2(_00909_),
    .B(_00916_),
    .C(_00912_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _16828_ (.A1(_03492_),
    .A2(_01821_),
    .A3(_00895_),
    .B1(_00893_),
    .B2(_00892_),
    .B3(_08464_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16829_ (.A1(_00890_),
    .A2(_00917_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16830_ (.I(_00918_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16831_ (.I(_00918_),
    .Z(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16832_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ),
    .A2(_00920_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16833_ (.I(_03509_),
    .Z(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16834_ (.A1(_01751_),
    .A2(_00919_),
    .B(_00921_),
    .C(_00922_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16835_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ),
    .A2(_00920_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16836_ (.A1(_01766_),
    .A2(_00919_),
    .B(_00923_),
    .C(_00922_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16837_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ),
    .A2(_00920_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16838_ (.A1(_08474_),
    .A2(_00919_),
    .B(_00924_),
    .C(_00922_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16839_ (.A1(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ),
    .A2(_00920_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16840_ (.A1(_00871_),
    .A2(_00919_),
    .B(_00925_),
    .C(_00922_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _16841_ (.A1(_08464_),
    .A2(_00860_),
    .A3(_00893_),
    .B1(_00906_),
    .B2(_01821_),
    .B3(_03492_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16842_ (.A1(_00890_),
    .A2(_00926_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16843_ (.I(_00927_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16844_ (.I(_00927_),
    .Z(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16845_ (.A1(_07822_),
    .A2(_00929_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16846_ (.I(_03509_),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16847_ (.A1(_01751_),
    .A2(_00928_),
    .B(_00930_),
    .C(_00931_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16848_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ),
    .A2(_00929_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16849_ (.A1(_01766_),
    .A2(_00928_),
    .B(_00932_),
    .C(_00931_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16850_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ),
    .A2(_00929_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16851_ (.A1(_01776_),
    .A2(_00928_),
    .B(_00933_),
    .C(_00931_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16852_ (.A1(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ),
    .A2(_00929_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16853_ (.A1(_00871_),
    .A2(_00928_),
    .B(_00934_),
    .C(_00931_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _16854_ (.A1(_03492_),
    .A2(_03496_),
    .A3(_00890_),
    .A4(_03525_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16855_ (.A1(\tt_um_rejunity_sn76489.noise[0].gen.restart_noise ),
    .A2(_04186_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16856_ (.A1(_00935_),
    .A2(_00936_),
    .B(_01828_),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16857_ (.I(\tt_um_rejunity_sn76489.latch_control_reg[0] ),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16858_ (.I(_03502_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16859_ (.I(_03766_),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16860_ (.A1(_03646_),
    .A2(_00938_),
    .B(_00939_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16861_ (.A1(_00937_),
    .A2(_00938_),
    .B(_00940_),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16862_ (.A1(_03493_),
    .A2(_03502_),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _16863_ (.A1(_00892_),
    .A2(_00938_),
    .B(_00941_),
    .C(_04129_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _16864_ (.A1(_00891_),
    .A2(_00938_),
    .B(_03526_),
    .C(_04129_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16865_ (.I(\tt_um_rejunity_sn76489.clk_counter[0] ),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16866_ (.A1(_00942_),
    .A2(_03759_),
    .B(_00939_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16867_ (.A1(_00942_),
    .A2(_03760_),
    .B(_00943_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16868_ (.A1(_00942_),
    .A2(_03759_),
    .B(\tt_um_rejunity_sn76489.clk_counter[1] ),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16869_ (.A1(\tt_um_rejunity_sn76489.clk_counter[1] ),
    .A2(_00942_),
    .A3(_03757_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _16870_ (.A1(_06941_),
    .A2(_00944_),
    .A3(_00945_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _16871_ (.A1(\tt_um_rejunity_sn76489.clk_counter[2] ),
    .A2(_00945_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16872_ (.A1(\tt_um_rejunity_sn76489.clk_counter[2] ),
    .A2(_00945_),
    .B(_01763_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16873_ (.A1(_00946_),
    .A2(_00947_),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16874_ (.A1(\tt_um_rejunity_sn76489.clk_counter[3] ),
    .A2(_00946_),
    .B(_00939_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16875_ (.A1(\tt_um_rejunity_sn76489.clk_counter[3] ),
    .A2(_00946_),
    .B(_00948_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16876_ (.A1(\tt_um_rejunity_sn76489.clk_counter[3] ),
    .A2(_00946_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _16877_ (.A1(\tt_um_rejunity_sn76489.clk_counter[4] ),
    .A2(_00949_),
    .Z(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16878_ (.A1(_08441_),
    .A2(_00950_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _16879_ (.A1(_01591_),
    .A2(_03756_),
    .B(_01052_),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16880_ (.I(_00951_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _16881_ (.I(_00951_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _16882_ (.A1(_01593_),
    .A2(_03764_),
    .B(_01103_),
    .C(_01080_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16883_ (.A1(_02709_),
    .A2(_03771_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16884_ (.A1(_03098_),
    .A2(_02754_),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _16885_ (.A1(_03545_),
    .A2(_03130_),
    .A3(_03133_),
    .A4(_00956_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _16886_ (.A1(_03775_),
    .A2(_00955_),
    .A3(_00957_),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _16887_ (.A1(_02709_),
    .A2(_03771_),
    .A3(_03130_),
    .A4(_02849_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _16888_ (.A1(_03797_),
    .A2(_03776_),
    .A3(_00956_),
    .A4(_00959_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16889_ (.A1(_00958_),
    .A2(_00960_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16890_ (.A1(_03774_),
    .A2(_03804_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _16891_ (.A1(_03797_),
    .A2(_03999_),
    .A3(_00955_),
    .A4(_00962_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _16892_ (.A1(_03774_),
    .A2(_03781_),
    .A3(_03804_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _16893_ (.A1(_03775_),
    .A2(_00955_),
    .A3(_00964_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _16894_ (.A1(_00961_),
    .A2(_00963_),
    .A3(_00965_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _16895_ (.A1(_01277_),
    .A2(_02457_),
    .B(\channels.clk_div[0] ),
    .C(_01105_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _16896_ (.A1(_03553_),
    .A2(_03784_),
    .A3(_00967_),
    .A4(_00966_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _16897_ (.I(_00968_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _16898_ (.I(_00969_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _16899_ (.A1(_00954_),
    .A2(_00966_),
    .B1(_00970_),
    .B2(_01193_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16900_ (.A1(_00953_),
    .A2(_00971_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16901_ (.A1(_01190_),
    .A2(_00952_),
    .B(_00972_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16902_ (.A1(_00955_),
    .A2(_00964_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16903_ (.A1(_03775_),
    .A2(_00973_),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16904_ (.A1(_00960_),
    .A2(_00974_),
    .B(_00954_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16905_ (.A1(_01221_),
    .A2(_00969_),
    .B(_00975_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16906_ (.A1(_00953_),
    .A2(_00976_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16907_ (.A1(_01218_),
    .A2(_00952_),
    .B(_00977_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _16908_ (.A1(_00954_),
    .A2(_00968_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16909_ (.A1(_01199_),
    .A2(_00970_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _16910_ (.A1(_00963_),
    .A2(_00978_),
    .B(_00979_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16911_ (.I0(_00980_),
    .I1(\channels.exp_periods[2][2] ),
    .S(_00951_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16912_ (.I(_00981_),
    .Z(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16913_ (.A1(_00958_),
    .A2(_00974_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _16914_ (.A1(_01215_),
    .A2(_00969_),
    .B1(_00978_),
    .B2(_00982_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16915_ (.A1(_00953_),
    .A2(_00983_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16916_ (.A1(_01212_),
    .A2(_00952_),
    .B(_00984_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _16917_ (.A1(_01206_),
    .A2(_00969_),
    .B1(_00973_),
    .B2(_00978_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _16918_ (.A1(_00953_),
    .A2(_00985_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16919_ (.A1(_01203_),
    .A2(_00952_),
    .B(_00986_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16920_ (.A1(_01593_),
    .A2(_03768_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _16921_ (.A1(_01826_),
    .A2(_00987_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16922_ (.I(_00988_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16923_ (.I0(_00971_),
    .I1(\channels.exp_periods[1][0] ),
    .S(_00989_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16924_ (.I(_00990_),
    .Z(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16925_ (.I0(_00976_),
    .I1(\channels.exp_periods[1][1] ),
    .S(_00989_),
    .Z(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16926_ (.I(_00991_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16927_ (.I0(_00980_),
    .I1(\channels.exp_periods[1][2] ),
    .S(_00989_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16928_ (.I(_00992_),
    .Z(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16929_ (.I0(_00983_),
    .I1(\channels.exp_periods[1][3] ),
    .S(_00989_),
    .Z(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16930_ (.I(_00993_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16931_ (.I0(_00985_),
    .I1(\channels.exp_periods[1][4] ),
    .S(_00988_),
    .Z(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16932_ (.I(_00994_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16933_ (.I(\channels.exp_counter[3][0] ),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16934_ (.I(_00995_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16935_ (.I(\channels.exp_counter[3][1] ),
    .Z(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16936_ (.I(_00996_),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16937_ (.I(\channels.exp_counter[3][2] ),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16938_ (.I(_00997_),
    .Z(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16939_ (.I(\channels.exp_counter[3][3] ),
    .Z(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16940_ (.I(_00998_),
    .Z(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16941_ (.I(\channels.exp_counter[3][4] ),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16942_ (.I(_00999_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _16943_ (.A1(_03773_),
    .A2(_03756_),
    .B(_01600_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16944_ (.I(_01000_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16945_ (.I0(_00971_),
    .I1(\channels.exp_periods[0][0] ),
    .S(_01001_),
    .Z(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16946_ (.I(_01002_),
    .Z(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16947_ (.I0(_00976_),
    .I1(\channels.exp_periods[0][1] ),
    .S(_01001_),
    .Z(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16948_ (.I(_01003_),
    .Z(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16949_ (.I0(_00980_),
    .I1(\channels.exp_periods[0][2] ),
    .S(_01001_),
    .Z(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16950_ (.I(_01004_),
    .Z(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16951_ (.I0(_00983_),
    .I1(\channels.exp_periods[0][3] ),
    .S(_01001_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16952_ (.I(_01005_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _16953_ (.I0(_00985_),
    .I1(\channels.exp_periods[0][4] ),
    .S(_01000_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _16954_ (.I(_01006_),
    .Z(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _16955_ (.A1(_01816_),
    .A2(_01810_),
    .A3(_03495_),
    .A4(_03502_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16956_ (.A1(\tt_um_rejunity_sn76489.control_noise[0][0] ),
    .A2(_01007_),
    .B(_00939_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16957_ (.A1(_01751_),
    .A2(_01007_),
    .B(_01008_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _16958_ (.A1(\tt_um_rejunity_sn76489.control_noise[0][1] ),
    .A2(_01007_),
    .B(_03767_),
    .ZN(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _16959_ (.A1(_08472_),
    .A2(_01007_),
    .B(_01009_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _16960_ (.A1(\tt_um_rejunity_sn76489.control_noise[0][2] ),
    .A2(_00935_),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _16961_ (.A1(_01776_),
    .A2(_00935_),
    .B(_01010_),
    .C(_07733_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16962_ (.D(_00011_),
    .CLK(clknet_leaf_190_clk),
    .Q(\channels.ring_outs[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16963_ (.D(_00012_),
    .CLK(clknet_leaf_190_clk),
    .Q(\channels.ring_outs[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16964_ (.D(_00013_),
    .CLK(clknet_leaf_212_clk),
    .Q(\channels.lfsr[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16965_ (.D(_00014_),
    .CLK(clknet_leaf_214_clk),
    .Q(\channels.lfsr[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16966_ (.D(_00015_),
    .CLK(clknet_leaf_213_clk),
    .Q(\channels.lfsr[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16967_ (.D(_00016_),
    .CLK(clknet_leaf_215_clk),
    .Q(\channels.lfsr[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16968_ (.D(_00017_),
    .CLK(clknet_leaf_219_clk),
    .Q(\channels.lfsr[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16969_ (.D(_00018_),
    .CLK(clknet_leaf_219_clk),
    .Q(\channels.lfsr[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16970_ (.D(_00019_),
    .CLK(clknet_leaf_219_clk),
    .Q(\channels.lfsr[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16971_ (.D(_00020_),
    .CLK(clknet_leaf_220_clk),
    .Q(\channels.lfsr[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16972_ (.D(_00021_),
    .CLK(clknet_leaf_221_clk),
    .Q(\channels.lfsr[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16973_ (.D(_00022_),
    .CLK(clknet_leaf_226_clk),
    .Q(\channels.lfsr[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16974_ (.D(_00023_),
    .CLK(clknet_leaf_226_clk),
    .Q(\channels.lfsr[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16975_ (.D(_00024_),
    .CLK(clknet_leaf_227_clk),
    .Q(\channels.lfsr[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16976_ (.D(_00025_),
    .CLK(clknet_leaf_227_clk),
    .Q(\channels.lfsr[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16977_ (.D(_00026_),
    .CLK(clknet_leaf_234_clk),
    .Q(\channels.lfsr[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16978_ (.D(_00027_),
    .CLK(clknet_leaf_235_clk),
    .Q(\channels.lfsr[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16979_ (.D(_00028_),
    .CLK(clknet_leaf_235_clk),
    .Q(\channels.lfsr[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16980_ (.D(_00029_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[3][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16981_ (.D(_00030_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16982_ (.D(_00031_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[3][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16983_ (.D(_00032_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16984_ (.D(_00033_),
    .CLK(clknet_leaf_230_clk),
    .Q(\channels.lfsr[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16985_ (.D(_00034_),
    .CLK(clknet_leaf_230_clk),
    .Q(\channels.lfsr[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16986_ (.D(_00035_),
    .CLK(clknet_leaf_210_clk),
    .Q(\channels.lfsr[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16987_ (.D(_00036_),
    .CLK(clknet_leaf_185_clk),
    .Q(\channels.env_vol[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16988_ (.D(_00037_),
    .CLK(clknet_leaf_185_clk),
    .Q(\channels.env_vol[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16989_ (.D(_00038_),
    .CLK(clknet_leaf_210_clk),
    .Q(\channels.env_vol[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16990_ (.D(_00039_),
    .CLK(clknet_leaf_209_clk),
    .Q(\channels.env_vol[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16991_ (.D(_00040_),
    .CLK(clknet_leaf_211_clk),
    .Q(\channels.env_vol[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16992_ (.D(_00041_),
    .CLK(clknet_leaf_209_clk),
    .Q(\channels.env_vol[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16993_ (.D(_00042_),
    .CLK(clknet_leaf_212_clk),
    .Q(\channels.env_vol[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16994_ (.D(_00043_),
    .CLK(clknet_leaf_209_clk),
    .Q(\channels.env_vol[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16995_ (.D(_00044_),
    .CLK(clknet_leaf_194_clk),
    .Q(\channels.exp_counter[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16996_ (.D(_00045_),
    .CLK(clknet_leaf_196_clk),
    .Q(\channels.exp_counter[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16997_ (.D(_00046_),
    .CLK(clknet_leaf_196_clk),
    .Q(\channels.exp_counter[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16998_ (.D(_00047_),
    .CLK(clknet_leaf_192_clk),
    .Q(\channels.exp_counter[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _16999_ (.D(_00048_),
    .CLK(clknet_leaf_192_clk),
    .Q(\channels.exp_counter[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17000_ (.D(_00049_),
    .CLK(clknet_leaf_194_clk),
    .Q(\channels.exp_counter[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17001_ (.D(_00050_),
    .CLK(clknet_leaf_194_clk),
    .Q(\channels.exp_counter[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17002_ (.D(_00051_),
    .CLK(clknet_5_23__leaf_clk),
    .Q(\channels.exp_counter[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17003_ (.D(_00052_),
    .CLK(clknet_leaf_193_clk),
    .Q(\channels.exp_counter[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17004_ (.D(_00053_),
    .CLK(clknet_leaf_191_clk),
    .Q(\channels.exp_counter[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17005_ (.D(_00054_),
    .CLK(clknet_leaf_194_clk),
    .Q(\channels.ring_outs[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17006_ (.D(_00055_),
    .CLK(clknet_leaf_183_clk),
    .Q(\channels.accum[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17007_ (.D(_00056_),
    .CLK(clknet_leaf_184_clk),
    .Q(\channels.accum[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17008_ (.D(_00057_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.accum[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17009_ (.D(_00058_),
    .CLK(clknet_5_18__leaf_clk),
    .Q(\channels.accum[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17010_ (.D(_00059_),
    .CLK(clknet_leaf_188_clk),
    .Q(\channels.accum[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17011_ (.D(_00060_),
    .CLK(clknet_leaf_172_clk),
    .Q(\channels.accum[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17012_ (.D(_00061_),
    .CLK(clknet_leaf_188_clk),
    .Q(\channels.accum[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17013_ (.D(_00062_),
    .CLK(clknet_leaf_171_clk),
    .Q(\channels.accum[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17014_ (.D(_00063_),
    .CLK(clknet_leaf_155_clk),
    .Q(\channels.accum[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17015_ (.D(_00064_),
    .CLK(clknet_leaf_167_clk),
    .Q(\channels.accum[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17016_ (.D(_00065_),
    .CLK(clknet_leaf_154_clk),
    .Q(\channels.accum[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17017_ (.D(_00066_),
    .CLK(clknet_leaf_150_clk),
    .Q(\channels.accum[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17018_ (.D(_00067_),
    .CLK(clknet_leaf_155_clk),
    .Q(\channels.accum[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17019_ (.D(_00068_),
    .CLK(clknet_leaf_150_clk),
    .Q(\channels.accum[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17020_ (.D(_00069_),
    .CLK(clknet_leaf_156_clk),
    .Q(\channels.accum[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17021_ (.D(_00070_),
    .CLK(clknet_leaf_163_clk),
    .Q(\channels.accum[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17022_ (.D(_00071_),
    .CLK(clknet_leaf_159_clk),
    .Q(\channels.accum[0][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17023_ (.D(_00072_),
    .CLK(clknet_leaf_193_clk),
    .Q(\channels.accum[0][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17024_ (.D(_00073_),
    .CLK(clknet_leaf_160_clk),
    .Q(\channels.accum[0][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17025_ (.D(_00074_),
    .CLK(clknet_leaf_162_clk),
    .Q(\channels.accum[0][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17026_ (.D(_00075_),
    .CLK(clknet_leaf_159_clk),
    .Q(\channels.accum[0][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17027_ (.D(_00076_),
    .CLK(clknet_leaf_193_clk),
    .Q(\channels.accum[0][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17028_ (.D(_00077_),
    .CLK(clknet_leaf_160_clk),
    .Q(\channels.accum[0][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17029_ (.D(_00078_),
    .CLK(clknet_leaf_161_clk),
    .Q(\channels.accum[0][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17030_ (.D(_00079_),
    .CLK(clknet_leaf_211_clk),
    .Q(\channels.lfsr[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17031_ (.D(_00080_),
    .CLK(clknet_leaf_210_clk),
    .Q(\channels.lfsr[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17032_ (.D(_00081_),
    .CLK(clknet_leaf_211_clk),
    .Q(\channels.lfsr[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17033_ (.D(_00082_),
    .CLK(clknet_leaf_217_clk),
    .Q(\channels.lfsr[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17034_ (.D(_00083_),
    .CLK(clknet_leaf_217_clk),
    .Q(\channels.lfsr[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17035_ (.D(_00084_),
    .CLK(clknet_leaf_223_clk),
    .Q(\channels.lfsr[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17036_ (.D(_00085_),
    .CLK(clknet_leaf_223_clk),
    .Q(\channels.lfsr[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17037_ (.D(_00086_),
    .CLK(clknet_leaf_222_clk),
    .Q(\channels.lfsr[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17038_ (.D(_00087_),
    .CLK(clknet_leaf_222_clk),
    .Q(\channels.lfsr[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17039_ (.D(_00088_),
    .CLK(clknet_leaf_225_clk),
    .Q(\channels.lfsr[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17040_ (.D(_00089_),
    .CLK(clknet_leaf_226_clk),
    .Q(\channels.lfsr[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17041_ (.D(_00090_),
    .CLK(clknet_leaf_227_clk),
    .Q(\channels.lfsr[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17042_ (.D(_00091_),
    .CLK(clknet_leaf_228_clk),
    .Q(\channels.lfsr[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17043_ (.D(_00092_),
    .CLK(clknet_leaf_234_clk),
    .Q(\channels.lfsr[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17044_ (.D(_00093_),
    .CLK(clknet_leaf_233_clk),
    .Q(\channels.lfsr[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17045_ (.D(_00094_),
    .CLK(clknet_leaf_235_clk),
    .Q(\channels.lfsr[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17046_ (.D(_00095_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17047_ (.D(_00096_),
    .CLK(clknet_leaf_233_clk),
    .Q(\channels.lfsr[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17048_ (.D(_00097_),
    .CLK(clknet_leaf_231_clk),
    .Q(\channels.lfsr[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17049_ (.D(_00098_),
    .CLK(clknet_leaf_232_clk),
    .Q(\channels.lfsr[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17050_ (.D(_00099_),
    .CLK(clknet_leaf_230_clk),
    .Q(\channels.lfsr[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17051_ (.D(_00100_),
    .CLK(clknet_leaf_230_clk),
    .Q(\channels.lfsr[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17052_ (.D(_00101_),
    .CLK(clknet_leaf_210_clk),
    .Q(\channels.lfsr[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17053_ (.D(_00000_),
    .CLK(clknet_leaf_90_clk),
    .Q(\filters.res_lut[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17054_ (.D(_00001_),
    .CLK(clknet_leaf_240_clk),
    .Q(\filters.res_lut[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17055_ (.D(_00002_),
    .CLK(clknet_leaf_91_clk),
    .Q(\filters.res_lut[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17056_ (.D(_00003_),
    .CLK(clknet_leaf_240_clk),
    .Q(\filters.res_lut[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17057_ (.D(_00004_),
    .CLK(clknet_leaf_90_clk),
    .Q(\filters.res_lut[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17058_ (.D(_00005_),
    .CLK(clknet_leaf_239_clk),
    .Q(\filters.res_lut[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17059_ (.D(_00006_),
    .CLK(clknet_leaf_84_clk),
    .Q(\filters.res_lut[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17060_ (.D(_00007_),
    .CLK(clknet_leaf_90_clk),
    .Q(\filters.res_lut[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17061_ (.D(_00008_),
    .CLK(clknet_leaf_85_clk),
    .Q(\filters.res_lut[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17062_ (.D(_00102_),
    .CLK(clknet_leaf_214_clk),
    .Q(\channels.lfsr[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17063_ (.D(_00103_),
    .CLK(clknet_leaf_215_clk),
    .Q(\channels.lfsr[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17064_ (.D(_00104_),
    .CLK(clknet_leaf_212_clk),
    .Q(\channels.lfsr[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17065_ (.D(_00105_),
    .CLK(clknet_leaf_216_clk),
    .Q(\channels.lfsr[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17066_ (.D(_00106_),
    .CLK(clknet_leaf_217_clk),
    .Q(\channels.lfsr[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17067_ (.D(_00107_),
    .CLK(clknet_leaf_218_clk),
    .Q(\channels.lfsr[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17068_ (.D(_00108_),
    .CLK(clknet_leaf_218_clk),
    .Q(\channels.lfsr[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17069_ (.D(_00109_),
    .CLK(clknet_leaf_221_clk),
    .Q(\channels.lfsr[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17070_ (.D(_00110_),
    .CLK(clknet_leaf_222_clk),
    .Q(\channels.lfsr[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17071_ (.D(_00111_),
    .CLK(clknet_leaf_224_clk),
    .Q(\channels.lfsr[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17072_ (.D(_00112_),
    .CLK(clknet_leaf_226_clk),
    .Q(\channels.lfsr[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17073_ (.D(_00113_),
    .CLK(clknet_leaf_225_clk),
    .Q(\channels.lfsr[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17074_ (.D(_00114_),
    .CLK(clknet_leaf_228_clk),
    .Q(\channels.lfsr[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17075_ (.D(_00115_),
    .CLK(clknet_leaf_234_clk),
    .Q(\channels.lfsr[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17076_ (.D(_00116_),
    .CLK(clknet_leaf_233_clk),
    .Q(\channels.lfsr[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17077_ (.D(_00117_),
    .CLK(clknet_leaf_235_clk),
    .Q(\channels.lfsr[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17078_ (.D(_00118_),
    .CLK(clknet_leaf_236_clk),
    .Q(\channels.lfsr[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17079_ (.D(_00119_),
    .CLK(clknet_leaf_233_clk),
    .Q(\channels.lfsr[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17080_ (.D(_00120_),
    .CLK(clknet_leaf_229_clk),
    .Q(\channels.lfsr[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17081_ (.D(_00121_),
    .CLK(clknet_leaf_232_clk),
    .Q(\channels.lfsr[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17082_ (.D(_00122_),
    .CLK(clknet_leaf_230_clk),
    .Q(\channels.lfsr[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17083_ (.D(_00123_),
    .CLK(clknet_leaf_224_clk),
    .Q(\channels.lfsr[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17084_ (.D(_00124_),
    .CLK(clknet_leaf_210_clk),
    .Q(\channels.lfsr[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17085_ (.D(_00125_),
    .CLK(clknet_leaf_89_clk),
    .Q(\filters.filt_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17086_ (.D(_00126_),
    .CLK(clknet_leaf_89_clk),
    .Q(\filters.filt_2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17087_ (.D(_00127_),
    .CLK(clknet_leaf_92_clk),
    .Q(\filters.filt_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17088_ (.D(_00128_),
    .CLK(clknet_leaf_74_clk),
    .Q(\filters.res_filt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17089_ (.D(_00129_),
    .CLK(clknet_leaf_86_clk),
    .Q(\filters.res_filt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17090_ (.D(_00130_),
    .CLK(clknet_leaf_86_clk),
    .Q(\filters.res_filt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17091_ (.D(_00131_),
    .CLK(clknet_leaf_88_clk),
    .Q(\filters.res_filt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17092_ (.D(_00132_),
    .CLK(clknet_leaf_87_clk),
    .Q(\filters.res_filt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17093_ (.D(_00133_),
    .CLK(clknet_leaf_74_clk),
    .Q(\filters.mode_vol[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17094_ (.D(_00134_),
    .CLK(clknet_5_15__leaf_clk),
    .Q(\filters.mode_vol[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17095_ (.D(_00135_),
    .CLK(clknet_leaf_108_clk),
    .Q(\filters.mode_vol[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17096_ (.D(_00136_),
    .CLK(clknet_leaf_108_clk),
    .Q(\filters.mode_vol[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17097_ (.D(_00137_),
    .CLK(clknet_leaf_69_clk),
    .Q(\filters.lp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17098_ (.D(_00138_),
    .CLK(clknet_leaf_69_clk),
    .Q(\filters.bp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17099_ (.D(_00139_),
    .CLK(clknet_leaf_69_clk),
    .Q(\filters.hp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17100_ (.D(_00140_),
    .CLK(clknet_leaf_69_clk),
    .Q(\filters.mode_vol[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17101_ (.D(_00141_),
    .CLK(clknet_leaf_105_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17102_ (.D(_00142_),
    .CLK(clknet_leaf_105_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17103_ (.D(_00143_),
    .CLK(clknet_leaf_115_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17104_ (.D(_00144_),
    .CLK(clknet_leaf_115_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17105_ (.D(_00145_),
    .CLK(clknet_leaf_121_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17106_ (.D(_00146_),
    .CLK(clknet_leaf_121_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17107_ (.D(_00147_),
    .CLK(clknet_leaf_121_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17108_ (.D(_00148_),
    .CLK(clknet_5_26__leaf_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17109_ (.D(_00149_),
    .CLK(clknet_leaf_109_clk),
    .Q(\channels.freq1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17110_ (.D(_00150_),
    .CLK(clknet_leaf_109_clk),
    .Q(\channels.freq1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17111_ (.D(_00151_),
    .CLK(clknet_leaf_109_clk),
    .Q(\channels.freq1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17112_ (.D(_00152_),
    .CLK(clknet_leaf_110_clk),
    .Q(\channels.freq1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17113_ (.D(_00153_),
    .CLK(clknet_leaf_109_clk),
    .Q(\channels.freq1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17114_ (.D(_00154_),
    .CLK(clknet_leaf_110_clk),
    .Q(\channels.freq1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17115_ (.D(_00155_),
    .CLK(clknet_leaf_110_clk),
    .Q(\channels.freq1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17116_ (.D(_00156_),
    .CLK(clknet_leaf_110_clk),
    .Q(\channels.freq1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17117_ (.D(_00157_),
    .CLK(clknet_leaf_108_clk),
    .Q(\channels.pw1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17118_ (.D(_00158_),
    .CLK(clknet_leaf_107_clk),
    .Q(\channels.pw1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17119_ (.D(_00159_),
    .CLK(clknet_leaf_107_clk),
    .Q(\channels.pw1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17120_ (.D(_00160_),
    .CLK(clknet_leaf_108_clk),
    .Q(\channels.pw1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17121_ (.D(_00161_),
    .CLK(clknet_leaf_113_clk),
    .Q(\channels.ctrl_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17122_ (.D(_00162_),
    .CLK(clknet_leaf_112_clk),
    .Q(\channels.ctrl_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17123_ (.D(_00163_),
    .CLK(clknet_leaf_112_clk),
    .Q(\channels.ctrl_reg1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17124_ (.D(_00164_),
    .CLK(clknet_leaf_113_clk),
    .Q(\channels.ctrl_reg1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17125_ (.D(_00165_),
    .CLK(clknet_leaf_112_clk),
    .Q(\channels.ctrl_reg1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17126_ (.D(_00166_),
    .CLK(clknet_leaf_68_clk),
    .Q(\channels.ctrl_reg1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17127_ (.D(_00167_),
    .CLK(clknet_leaf_68_clk),
    .Q(\channels.ctrl_reg1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17128_ (.D(_00168_),
    .CLK(clknet_leaf_68_clk),
    .Q(\channels.ctrl_reg1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17129_ (.D(_00169_),
    .CLK(clknet_leaf_114_clk),
    .Q(\channels.atk_dec1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17130_ (.D(_00170_),
    .CLK(clknet_leaf_114_clk),
    .Q(\channels.atk_dec1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17131_ (.D(_00171_),
    .CLK(clknet_leaf_114_clk),
    .Q(\channels.atk_dec1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17132_ (.D(_00172_),
    .CLK(clknet_leaf_114_clk),
    .Q(\channels.atk_dec1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17133_ (.D(_00173_),
    .CLK(clknet_leaf_111_clk),
    .Q(\channels.atk_dec1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17134_ (.D(_00174_),
    .CLK(clknet_leaf_112_clk),
    .Q(\channels.atk_dec1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17135_ (.D(_00175_),
    .CLK(clknet_leaf_111_clk),
    .Q(\channels.atk_dec1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17136_ (.D(_00176_),
    .CLK(clknet_leaf_111_clk),
    .Q(\channels.atk_dec1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17137_ (.D(_00177_),
    .CLK(clknet_leaf_114_clk),
    .Q(\channels.sus_rel1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17138_ (.D(_00178_),
    .CLK(clknet_leaf_113_clk),
    .Q(\channels.sus_rel1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17139_ (.D(_00179_),
    .CLK(clknet_leaf_113_clk),
    .Q(\channels.sus_rel1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17140_ (.D(_00180_),
    .CLK(clknet_leaf_113_clk),
    .Q(\channels.sus_rel1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17141_ (.D(_00181_),
    .CLK(clknet_leaf_117_clk),
    .Q(\channels.sus_rel1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17142_ (.D(_00182_),
    .CLK(clknet_leaf_117_clk),
    .Q(\channels.sus_rel1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17143_ (.D(_00183_),
    .CLK(clknet_leaf_117_clk),
    .Q(\channels.sus_rel1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17144_ (.D(_00184_),
    .CLK(clknet_leaf_117_clk),
    .Q(\channels.sus_rel1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17145_ (.D(_00185_),
    .CLK(clknet_leaf_116_clk),
    .Q(\channels.freq2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17146_ (.D(_00186_),
    .CLK(clknet_leaf_114_clk),
    .Q(\channels.freq2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17147_ (.D(_00187_),
    .CLK(clknet_leaf_114_clk),
    .Q(\channels.freq2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17148_ (.D(_00188_),
    .CLK(clknet_leaf_115_clk),
    .Q(\channels.freq2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17149_ (.D(_00189_),
    .CLK(clknet_leaf_115_clk),
    .Q(\channels.freq2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17150_ (.D(_00190_),
    .CLK(clknet_leaf_116_clk),
    .Q(\channels.freq2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17151_ (.D(_00191_),
    .CLK(clknet_leaf_118_clk),
    .Q(\channels.freq2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17152_ (.D(_00192_),
    .CLK(clknet_leaf_118_clk),
    .Q(\channels.freq2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17153_ (.D(_00193_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.pw2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17154_ (.D(_00194_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.pw2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17155_ (.D(_00195_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.pw2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17156_ (.D(_00196_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.pw2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17157_ (.D(_00197_),
    .CLK(clknet_leaf_128_clk),
    .Q(\channels.ctrl_reg2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17158_ (.D(_00198_),
    .CLK(clknet_leaf_128_clk),
    .Q(\channels.ctrl_reg2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17159_ (.D(_00199_),
    .CLK(clknet_leaf_128_clk),
    .Q(\channels.ctrl_reg2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17160_ (.D(_00200_),
    .CLK(clknet_leaf_119_clk),
    .Q(\channels.ctrl_reg2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17161_ (.D(_00201_),
    .CLK(clknet_leaf_119_clk),
    .Q(\channels.ctrl_reg2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17162_ (.D(_00202_),
    .CLK(clknet_leaf_118_clk),
    .Q(\channels.ctrl_reg2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17163_ (.D(_00203_),
    .CLK(clknet_leaf_118_clk),
    .Q(\channels.ctrl_reg2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17164_ (.D(_00204_),
    .CLK(clknet_leaf_119_clk),
    .Q(\channels.ctrl_reg2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17165_ (.D(_00205_),
    .CLK(clknet_leaf_127_clk),
    .Q(\channels.atk_dec2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17166_ (.D(_00206_),
    .CLK(clknet_leaf_126_clk),
    .Q(\channels.atk_dec2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17167_ (.D(_00207_),
    .CLK(clknet_leaf_126_clk),
    .Q(\channels.atk_dec2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17168_ (.D(_00208_),
    .CLK(clknet_leaf_126_clk),
    .Q(\channels.atk_dec2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17169_ (.D(_00209_),
    .CLK(clknet_leaf_120_clk),
    .Q(\channels.atk_dec2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17170_ (.D(_00210_),
    .CLK(clknet_leaf_120_clk),
    .Q(\channels.atk_dec2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17171_ (.D(_00211_),
    .CLK(clknet_leaf_120_clk),
    .Q(\channels.atk_dec2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17172_ (.D(_00212_),
    .CLK(clknet_leaf_120_clk),
    .Q(\channels.atk_dec2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17173_ (.D(_00213_),
    .CLK(clknet_leaf_127_clk),
    .Q(\channels.sus_rel2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17174_ (.D(_00214_),
    .CLK(clknet_leaf_125_clk),
    .Q(\channels.sus_rel2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17175_ (.D(_00215_),
    .CLK(clknet_leaf_125_clk),
    .Q(\channels.sus_rel2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17176_ (.D(_00216_),
    .CLK(clknet_leaf_131_clk),
    .Q(\channels.sus_rel2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17177_ (.D(_00217_),
    .CLK(clknet_leaf_147_clk),
    .Q(\channels.sus_rel2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17178_ (.D(_00218_),
    .CLK(clknet_leaf_147_clk),
    .Q(\channels.sus_rel2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17179_ (.D(_00219_),
    .CLK(clknet_leaf_146_clk),
    .Q(\channels.sus_rel2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17180_ (.D(_00220_),
    .CLK(clknet_leaf_146_clk),
    .Q(\channels.sus_rel2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17181_ (.D(_00221_),
    .CLK(clknet_leaf_144_clk),
    .Q(\channels.freq3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17182_ (.D(_00222_),
    .CLK(clknet_leaf_144_clk),
    .Q(\channels.freq3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17183_ (.D(_00223_),
    .CLK(clknet_leaf_144_clk),
    .Q(\channels.freq3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17184_ (.D(_00224_),
    .CLK(clknet_leaf_144_clk),
    .Q(\channels.freq3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17185_ (.D(_00225_),
    .CLK(clknet_leaf_123_clk),
    .Q(\channels.freq3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17186_ (.D(_00226_),
    .CLK(clknet_leaf_123_clk),
    .Q(\channels.freq3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17187_ (.D(_00227_),
    .CLK(clknet_leaf_146_clk),
    .Q(\channels.freq3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17188_ (.D(_00228_),
    .CLK(clknet_leaf_123_clk),
    .Q(\channels.freq3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17189_ (.D(_00229_),
    .CLK(clknet_leaf_145_clk),
    .Q(\channels.pw3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17190_ (.D(_00230_),
    .CLK(clknet_leaf_145_clk),
    .Q(\channels.pw3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17191_ (.D(_00231_),
    .CLK(clknet_leaf_145_clk),
    .Q(\channels.pw3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17192_ (.D(_00232_),
    .CLK(clknet_leaf_143_clk),
    .Q(\channels.pw3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17193_ (.D(_00233_),
    .CLK(clknet_leaf_152_clk),
    .Q(\channels.ctrl_reg3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17194_ (.D(_00234_),
    .CLK(clknet_leaf_148_clk),
    .Q(\channels.ctrl_reg3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17195_ (.D(_00235_),
    .CLK(clknet_leaf_149_clk),
    .Q(\channels.ctrl_reg3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17196_ (.D(_00236_),
    .CLK(clknet_leaf_145_clk),
    .Q(\channels.ctrl_reg3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17197_ (.D(_00237_),
    .CLK(clknet_leaf_148_clk),
    .Q(\channels.ctrl_reg3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17198_ (.D(_00238_),
    .CLK(clknet_leaf_168_clk),
    .Q(\channels.ctrl_reg3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17199_ (.D(_00239_),
    .CLK(clknet_leaf_148_clk),
    .Q(\channels.ctrl_reg3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17200_ (.D(_00240_),
    .CLK(clknet_leaf_168_clk),
    .Q(\channels.ctrl_reg3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17201_ (.D(_00241_),
    .CLK(clknet_leaf_124_clk),
    .Q(\channels.atk_dec3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17202_ (.D(_00242_),
    .CLK(clknet_leaf_125_clk),
    .Q(\channels.atk_dec3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17203_ (.D(_00243_),
    .CLK(clknet_leaf_144_clk),
    .Q(\channels.atk_dec3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17204_ (.D(_00244_),
    .CLK(clknet_leaf_125_clk),
    .Q(\channels.atk_dec3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17205_ (.D(_00245_),
    .CLK(clknet_leaf_124_clk),
    .Q(\channels.atk_dec3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17206_ (.D(_00246_),
    .CLK(clknet_leaf_124_clk),
    .Q(\channels.atk_dec3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17207_ (.D(_00247_),
    .CLK(clknet_leaf_124_clk),
    .Q(\channels.atk_dec3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17208_ (.D(_00248_),
    .CLK(clknet_leaf_126_clk),
    .Q(\channels.atk_dec3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17209_ (.D(_00249_),
    .CLK(clknet_leaf_74_clk),
    .Q(\channels.sus_rel3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17210_ (.D(_00250_),
    .CLK(clknet_leaf_73_clk),
    .Q(\channels.sus_rel3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17211_ (.D(_00251_),
    .CLK(clknet_leaf_73_clk),
    .Q(\channels.sus_rel3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17212_ (.D(_00252_),
    .CLK(clknet_leaf_73_clk),
    .Q(\channels.sus_rel3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17213_ (.D(_00253_),
    .CLK(clknet_leaf_76_clk),
    .Q(\channels.sus_rel3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17214_ (.D(_00254_),
    .CLK(clknet_leaf_86_clk),
    .Q(\channels.sus_rel3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17215_ (.D(_00255_),
    .CLK(clknet_leaf_75_clk),
    .Q(\channels.sus_rel3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17216_ (.D(_00256_),
    .CLK(clknet_leaf_75_clk),
    .Q(\channels.sus_rel3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17217_ (.D(_00257_),
    .CLK(clknet_leaf_77_clk),
    .Q(\filters.cutoff_lut[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17218_ (.D(_00258_),
    .CLK(clknet_leaf_78_clk),
    .Q(\filters.cutoff_lut[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17219_ (.D(_00259_),
    .CLK(clknet_leaf_73_clk),
    .Q(\filters.cutoff_lut[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17220_ (.D(_00260_),
    .CLK(clknet_leaf_78_clk),
    .Q(\filters.cutoff_lut[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17221_ (.D(_00261_),
    .CLK(clknet_leaf_76_clk),
    .Q(\filters.cutoff_lut[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17222_ (.D(_00262_),
    .CLK(clknet_leaf_86_clk),
    .Q(\filters.cutoff_lut[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17223_ (.D(_00263_),
    .CLK(clknet_leaf_77_clk),
    .Q(\filters.cutoff_lut[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17224_ (.D(_00264_),
    .CLK(clknet_leaf_77_clk),
    .Q(\filters.cutoff_lut[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17225_ (.D(_00265_),
    .CLK(clknet_leaf_47_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.signal_edge.previous_signal_state_0 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17226_ (.D(_00266_),
    .CLK(clknet_leaf_77_clk),
    .Q(\clk_trg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17227_ (.D(_00267_),
    .CLK(clknet_leaf_80_clk),
    .Q(\clk_trg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17228_ (.D(_00268_),
    .CLK(clknet_leaf_171_clk),
    .Q(\channels.sync_outs[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17229_ (.D(_00269_),
    .CLK(clknet_leaf_165_clk),
    .Q(\channels.sync_outs[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17230_ (.D(_00270_),
    .CLK(clknet_leaf_165_clk),
    .Q(\channels.sync_outs[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17231_ (.D(_00271_),
    .CLK(clknet_leaf_181_clk),
    .Q(\channels.sample3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17232_ (.D(_00272_),
    .CLK(clknet_leaf_180_clk),
    .Q(\channels.sample3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17233_ (.D(_00273_),
    .CLK(clknet_leaf_180_clk),
    .Q(\channels.sample3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17234_ (.D(_00274_),
    .CLK(clknet_leaf_178_clk),
    .Q(\channels.sample3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17235_ (.D(_00275_),
    .CLK(clknet_leaf_178_clk),
    .Q(\channels.sample3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17236_ (.D(_00276_),
    .CLK(clknet_leaf_177_clk),
    .Q(\channels.sample3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17237_ (.D(_00277_),
    .CLK(clknet_leaf_176_clk),
    .Q(\channels.sample3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17238_ (.D(_00278_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\channels.sample3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17239_ (.D(_00279_),
    .CLK(clknet_leaf_175_clk),
    .Q(\channels.sample3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17240_ (.D(_00280_),
    .CLK(clknet_leaf_95_clk),
    .Q(\channels.sample3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17241_ (.D(_00281_),
    .CLK(clknet_leaf_175_clk),
    .Q(\channels.sample3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17242_ (.D(_00282_),
    .CLK(clknet_leaf_174_clk),
    .Q(\channels.sample3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17243_ (.D(_00283_),
    .CLK(clknet_leaf_181_clk),
    .Q(\channels.sample2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17244_ (.D(_00284_),
    .CLK(clknet_leaf_180_clk),
    .Q(\channels.sample2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17245_ (.D(_00285_),
    .CLK(clknet_leaf_179_clk),
    .Q(\channels.sample2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17246_ (.D(_00286_),
    .CLK(clknet_leaf_178_clk),
    .Q(\channels.sample2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17247_ (.D(_00287_),
    .CLK(clknet_leaf_177_clk),
    .Q(\channels.sample2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17248_ (.D(_00288_),
    .CLK(clknet_leaf_177_clk),
    .Q(\channels.sample2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17249_ (.D(_00289_),
    .CLK(clknet_leaf_177_clk),
    .Q(\channels.sample2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17250_ (.D(_00290_),
    .CLK(clknet_leaf_176_clk),
    .Q(\channels.sample2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17251_ (.D(_00291_),
    .CLK(clknet_leaf_176_clk),
    .Q(\channels.sample2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17252_ (.D(_00292_),
    .CLK(clknet_leaf_96_clk),
    .Q(\channels.sample2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17253_ (.D(_00293_),
    .CLK(clknet_leaf_96_clk),
    .Q(\channels.sample2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17254_ (.D(_00294_),
    .CLK(clknet_leaf_174_clk),
    .Q(\channels.sample2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17255_ (.D(_00295_),
    .CLK(clknet_leaf_173_clk),
    .Q(\channels.sample1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17256_ (.D(_00296_),
    .CLK(clknet_leaf_178_clk),
    .Q(\channels.sample1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17257_ (.D(_00297_),
    .CLK(clknet_leaf_178_clk),
    .Q(\channels.sample1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17258_ (.D(_00298_),
    .CLK(clknet_leaf_181_clk),
    .Q(\channels.sample1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17259_ (.D(_00299_),
    .CLK(clknet_leaf_181_clk),
    .Q(\channels.sample1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17260_ (.D(_00300_),
    .CLK(clknet_leaf_177_clk),
    .Q(\channels.sample1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17261_ (.D(_00301_),
    .CLK(clknet_leaf_173_clk),
    .Q(\channels.sample1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17262_ (.D(_00302_),
    .CLK(clknet_leaf_176_clk),
    .Q(\channels.sample1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17263_ (.D(_00303_),
    .CLK(clknet_leaf_174_clk),
    .Q(\channels.sample1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17264_ (.D(_00304_),
    .CLK(clknet_leaf_175_clk),
    .Q(\channels.sample1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17265_ (.D(_00305_),
    .CLK(clknet_leaf_175_clk),
    .Q(\channels.sample1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17266_ (.D(_00306_),
    .CLK(clknet_leaf_174_clk),
    .Q(\channels.sample1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17267_ (.D(_00307_),
    .CLK(clknet_leaf_11_clk),
    .Q(\filters.sample_filtered[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17268_ (.D(_00308_),
    .CLK(clknet_leaf_11_clk),
    .Q(\filters.sample_filtered[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17269_ (.D(_00309_),
    .CLK(clknet_leaf_7_clk),
    .Q(\filters.sample_filtered[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17270_ (.D(_00310_),
    .CLK(clknet_leaf_9_clk),
    .Q(\filters.sample_filtered[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17271_ (.D(_00311_),
    .CLK(clknet_leaf_9_clk),
    .Q(\filters.sample_filtered[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17272_ (.D(_00312_),
    .CLK(clknet_leaf_10_clk),
    .Q(\filters.sample_filtered[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17273_ (.D(_00313_),
    .CLK(clknet_leaf_10_clk),
    .Q(\filters.sample_filtered[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17274_ (.D(_00314_),
    .CLK(clknet_5_7__leaf_clk),
    .Q(\filters.sample_filtered[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17275_ (.D(_00315_),
    .CLK(clknet_leaf_92_clk),
    .Q(\filters.sample_filtered[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17276_ (.D(_00316_),
    .CLK(clknet_leaf_91_clk),
    .Q(\filters.sample_filtered[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17277_ (.D(_00317_),
    .CLK(clknet_leaf_90_clk),
    .Q(\filters.sample_filtered[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17278_ (.D(_00318_),
    .CLK(clknet_leaf_90_clk),
    .Q(\filters.sample_filtered[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17279_ (.D(_00319_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\filters.sample_filtered[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17280_ (.D(_00320_),
    .CLK(clknet_leaf_14_clk),
    .Q(\filters.sample_filtered[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17281_ (.D(_00321_),
    .CLK(clknet_leaf_84_clk),
    .Q(\filters.sample_filtered[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17282_ (.D(_00322_),
    .CLK(clknet_leaf_17_clk),
    .Q(\filters.sample_filtered[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17283_ (.D(_00323_),
    .CLK(clknet_leaf_77_clk),
    .Q(\filters.cutoff_lut[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17284_ (.D(_00324_),
    .CLK(clknet_leaf_72_clk),
    .Q(\filters.cutoff_lut[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17285_ (.D(_00325_),
    .CLK(clknet_leaf_72_clk),
    .Q(\filters.cutoff_lut[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17286_ (.D(_00326_),
    .CLK(clknet_leaf_67_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17287_ (.D(_00327_),
    .CLK(clknet_leaf_71_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17288_ (.D(_00328_),
    .CLK(clknet_leaf_69_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17289_ (.D(_00329_),
    .CLK(clknet_leaf_67_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17290_ (.D(_00330_),
    .CLK(clknet_leaf_66_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17291_ (.D(_00331_),
    .CLK(clknet_leaf_67_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17292_ (.D(_00332_),
    .CLK(clknet_leaf_67_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17293_ (.D(_00333_),
    .CLK(clknet_leaf_66_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17294_ (.D(_00334_),
    .CLK(clknet_leaf_67_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17295_ (.D(_00335_),
    .CLK(clknet_leaf_67_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17296_ (.D(_00336_),
    .CLK(clknet_leaf_68_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17297_ (.D(_00337_),
    .CLK(clknet_leaf_69_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17298_ (.D(_00338_),
    .CLK(clknet_leaf_165_clk),
    .Q(\channels.adsr_state[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17299_ (.D(_00339_),
    .CLK(clknet_leaf_166_clk),
    .Q(\channels.adsr_state[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17300_ (.D(_00340_),
    .CLK(clknet_leaf_187_clk),
    .Q(\channels.accum[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17301_ (.D(_00341_),
    .CLK(clknet_leaf_184_clk),
    .Q(\channels.accum[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17302_ (.D(_00342_),
    .CLK(clknet_leaf_187_clk),
    .Q(\channels.accum[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17303_ (.D(_00343_),
    .CLK(clknet_leaf_180_clk),
    .Q(\channels.accum[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17304_ (.D(_00344_),
    .CLK(clknet_leaf_183_clk),
    .Q(\channels.accum[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17305_ (.D(_00345_),
    .CLK(clknet_leaf_173_clk),
    .Q(\channels.accum[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17306_ (.D(_00346_),
    .CLK(clknet_leaf_183_clk),
    .Q(\channels.accum[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17307_ (.D(_00347_),
    .CLK(clknet_leaf_172_clk),
    .Q(\channels.accum[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17308_ (.D(_00348_),
    .CLK(clknet_leaf_157_clk),
    .Q(\channels.accum[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17309_ (.D(_00349_),
    .CLK(clknet_leaf_167_clk),
    .Q(\channels.accum[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17310_ (.D(_00350_),
    .CLK(clknet_leaf_151_clk),
    .Q(\channels.accum[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17311_ (.D(_00351_),
    .CLK(clknet_leaf_149_clk),
    .Q(\channels.accum[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17312_ (.D(_00352_),
    .CLK(clknet_leaf_157_clk),
    .Q(\channels.accum[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17313_ (.D(_00353_),
    .CLK(clknet_leaf_166_clk),
    .Q(\channels.accum[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17314_ (.D(_00354_),
    .CLK(clknet_leaf_157_clk),
    .Q(\channels.accum[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17315_ (.D(_00355_),
    .CLK(clknet_leaf_163_clk),
    .Q(\channels.accum[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17316_ (.D(_00356_),
    .CLK(clknet_leaf_162_clk),
    .Q(\channels.accum[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17317_ (.D(_00357_),
    .CLK(clknet_leaf_190_clk),
    .Q(\channels.accum[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17318_ (.D(_00358_),
    .CLK(clknet_leaf_161_clk),
    .Q(\channels.accum[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17319_ (.D(_00359_),
    .CLK(clknet_leaf_163_clk),
    .Q(\channels.accum[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17320_ (.D(_00360_),
    .CLK(clknet_leaf_162_clk),
    .Q(\channels.accum[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17321_ (.D(_00361_),
    .CLK(clknet_leaf_190_clk),
    .Q(\channels.accum[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17322_ (.D(_00362_),
    .CLK(clknet_leaf_162_clk),
    .Q(\channels.accum[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17323_ (.D(_00363_),
    .CLK(clknet_leaf_164_clk),
    .Q(\channels.accum[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17324_ (.D(_00364_),
    .CLK(clknet_leaf_187_clk),
    .Q(\channels.accum[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17325_ (.D(_00365_),
    .CLK(clknet_leaf_184_clk),
    .Q(\channels.accum[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17326_ (.D(_00366_),
    .CLK(clknet_5_19__leaf_clk),
    .Q(\channels.accum[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17327_ (.D(_00367_),
    .CLK(clknet_leaf_180_clk),
    .Q(\channels.accum[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17328_ (.D(_00368_),
    .CLK(clknet_leaf_187_clk),
    .Q(\channels.accum[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17329_ (.D(_00369_),
    .CLK(clknet_leaf_181_clk),
    .Q(\channels.accum[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17330_ (.D(_00370_),
    .CLK(clknet_leaf_188_clk),
    .Q(\channels.accum[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17331_ (.D(_00371_),
    .CLK(clknet_leaf_172_clk),
    .Q(\channels.accum[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17332_ (.D(_00372_),
    .CLK(clknet_leaf_156_clk),
    .Q(\channels.accum[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17333_ (.D(_00373_),
    .CLK(clknet_leaf_150_clk),
    .Q(\channels.accum[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17334_ (.D(_00374_),
    .CLK(clknet_leaf_154_clk),
    .Q(\channels.accum[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17335_ (.D(_00375_),
    .CLK(clknet_leaf_149_clk),
    .Q(\channels.accum[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17336_ (.D(_00376_),
    .CLK(clknet_leaf_155_clk),
    .Q(\channels.accum[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17337_ (.D(_00377_),
    .CLK(clknet_leaf_167_clk),
    .Q(\channels.accum[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17338_ (.D(_00378_),
    .CLK(clknet_leaf_156_clk),
    .Q(\channels.accum[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17339_ (.D(_00379_),
    .CLK(clknet_leaf_163_clk),
    .Q(\channels.accum[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17340_ (.D(_00380_),
    .CLK(clknet_leaf_159_clk),
    .Q(\channels.accum[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17341_ (.D(_00381_),
    .CLK(clknet_leaf_190_clk),
    .Q(\channels.accum[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17342_ (.D(_00382_),
    .CLK(clknet_leaf_161_clk),
    .Q(\channels.accum[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17343_ (.D(_00383_),
    .CLK(clknet_leaf_163_clk),
    .Q(\channels.accum[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17344_ (.D(_00384_),
    .CLK(clknet_leaf_158_clk),
    .Q(\channels.accum[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17345_ (.D(_00385_),
    .CLK(clknet_leaf_190_clk),
    .Q(\channels.accum[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17346_ (.D(_00386_),
    .CLK(clknet_leaf_160_clk),
    .Q(\channels.accum[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17347_ (.D(_00387_),
    .CLK(clknet_leaf_164_clk),
    .Q(\channels.accum[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17348_ (.D(_00388_),
    .CLK(clknet_leaf_85_clk),
    .Q(\filters.res_lut[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17349_ (.D(_00389_),
    .CLK(clknet_leaf_85_clk),
    .Q(\filters.res_lut[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17350_ (.D(_00390_),
    .CLK(clknet_leaf_75_clk),
    .Q(\channels.freq1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17351_ (.D(_00391_),
    .CLK(clknet_leaf_75_clk),
    .Q(\channels.freq1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17352_ (.D(_00392_),
    .CLK(clknet_leaf_107_clk),
    .Q(\channels.freq1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17353_ (.D(_00393_),
    .CLK(clknet_leaf_107_clk),
    .Q(\channels.freq1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17354_ (.D(_00394_),
    .CLK(clknet_leaf_102_clk),
    .Q(\channels.freq1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17355_ (.D(_00395_),
    .CLK(clknet_leaf_101_clk),
    .Q(\channels.freq1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17356_ (.D(_00396_),
    .CLK(clknet_leaf_87_clk),
    .Q(\channels.freq1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17357_ (.D(_00397_),
    .CLK(clknet_leaf_75_clk),
    .Q(\channels.freq1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17358_ (.D(_00398_),
    .CLK(clknet_leaf_88_clk),
    .Q(\channels.pw1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17359_ (.D(_00399_),
    .CLK(clknet_leaf_87_clk),
    .Q(\channels.pw1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17360_ (.D(_00400_),
    .CLK(clknet_leaf_100_clk),
    .Q(\channels.pw1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17361_ (.D(_00401_),
    .CLK(clknet_leaf_99_clk),
    .Q(\channels.pw1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17362_ (.D(_00402_),
    .CLK(clknet_leaf_103_clk),
    .Q(\channels.pw1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17363_ (.D(_00403_),
    .CLK(clknet_leaf_87_clk),
    .Q(\channels.pw1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17364_ (.D(_00404_),
    .CLK(clknet_leaf_88_clk),
    .Q(\channels.pw1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17365_ (.D(_00405_),
    .CLK(clknet_leaf_99_clk),
    .Q(\channels.pw1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17366_ (.D(_00406_),
    .CLK(clknet_leaf_101_clk),
    .Q(\channels.freq2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17367_ (.D(_00407_),
    .CLK(clknet_leaf_101_clk),
    .Q(\channels.freq2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17368_ (.D(_00408_),
    .CLK(clknet_leaf_107_clk),
    .Q(\channels.freq2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17369_ (.D(_00409_),
    .CLK(clknet_leaf_106_clk),
    .Q(\channels.freq2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17370_ (.D(_00410_),
    .CLK(clknet_leaf_102_clk),
    .Q(\channels.freq2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17371_ (.D(_00411_),
    .CLK(clknet_leaf_102_clk),
    .Q(\channels.freq2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17372_ (.D(_00412_),
    .CLK(clknet_leaf_106_clk),
    .Q(\channels.freq2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17373_ (.D(_00413_),
    .CLK(clknet_leaf_106_clk),
    .Q(\channels.freq2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17374_ (.D(_00414_),
    .CLK(clknet_leaf_98_clk),
    .Q(\channels.freq3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17375_ (.D(_00415_),
    .CLK(clknet_leaf_100_clk),
    .Q(\channels.freq3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17376_ (.D(_00416_),
    .CLK(clknet_leaf_102_clk),
    .Q(\channels.freq3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17377_ (.D(_00417_),
    .CLK(clknet_leaf_99_clk),
    .Q(\channels.freq3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17378_ (.D(_00418_),
    .CLK(clknet_5_24__leaf_clk),
    .Q(\channels.freq3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17379_ (.D(_00419_),
    .CLK(clknet_leaf_103_clk),
    .Q(\channels.freq3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17380_ (.D(_00420_),
    .CLK(clknet_leaf_103_clk),
    .Q(\channels.freq3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17381_ (.D(_00421_),
    .CLK(clknet_leaf_103_clk),
    .Q(\channels.freq3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17382_ (.D(_00422_),
    .CLK(clknet_leaf_98_clk),
    .Q(\channels.pw3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17383_ (.D(_00423_),
    .CLK(clknet_leaf_98_clk),
    .Q(\channels.pw3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17384_ (.D(_00424_),
    .CLK(clknet_leaf_96_clk),
    .Q(\channels.pw3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17385_ (.D(_00425_),
    .CLK(clknet_leaf_95_clk),
    .Q(\channels.pw3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17386_ (.D(_00426_),
    .CLK(clknet_leaf_103_clk),
    .Q(\channels.pw3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17387_ (.D(_00427_),
    .CLK(clknet_leaf_97_clk),
    .Q(\channels.pw3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17388_ (.D(_00428_),
    .CLK(clknet_leaf_103_clk),
    .Q(\channels.pw3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17389_ (.D(_00429_),
    .CLK(clknet_leaf_97_clk),
    .Q(\channels.pw3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17390_ (.D(_00430_),
    .CLK(clknet_leaf_99_clk),
    .Q(\channels.pw2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17391_ (.D(_00431_),
    .CLK(clknet_leaf_98_clk),
    .Q(\channels.pw2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17392_ (.D(_00432_),
    .CLK(clknet_leaf_95_clk),
    .Q(\channels.pw2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17393_ (.D(_00433_),
    .CLK(clknet_leaf_95_clk),
    .Q(\channels.pw2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17394_ (.D(_00434_),
    .CLK(clknet_leaf_88_clk),
    .Q(\channels.pw2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17395_ (.D(_00435_),
    .CLK(clknet_leaf_99_clk),
    .Q(\channels.pw2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17396_ (.D(_00436_),
    .CLK(clknet_leaf_88_clk),
    .Q(\channels.pw2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17397_ (.D(_00437_),
    .CLK(clknet_leaf_88_clk),
    .Q(\channels.pw2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17398_ (.D(_00438_),
    .CLK(clknet_leaf_175_clk),
    .Q(\channels.clk_div[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17399_ (.D(_00439_),
    .CLK(clknet_leaf_169_clk),
    .Q(\channels.clk_div[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17400_ (.D(_00440_),
    .CLK(clknet_leaf_169_clk),
    .Q(\channels.clk_div[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17401_ (.D(_00441_),
    .CLK(clknet_leaf_207_clk),
    .Q(\channels.env_vol[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17402_ (.D(_00442_),
    .CLK(clknet_leaf_208_clk),
    .Q(\channels.env_vol[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17403_ (.D(_00443_),
    .CLK(clknet_leaf_207_clk),
    .Q(\channels.env_vol[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17404_ (.D(_00444_),
    .CLK(clknet_leaf_207_clk),
    .Q(\channels.env_vol[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17405_ (.D(_00445_),
    .CLK(clknet_leaf_211_clk),
    .Q(\channels.env_vol[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17406_ (.D(_00446_),
    .CLK(clknet_leaf_207_clk),
    .Q(\channels.env_vol[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17407_ (.D(_00447_),
    .CLK(clknet_leaf_204_clk),
    .Q(\channels.env_vol[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17408_ (.D(_00448_),
    .CLK(clknet_leaf_204_clk),
    .Q(\channels.env_vol[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17409_ (.D(_00449_),
    .CLK(clknet_leaf_132_clk),
    .Q(\channels.env_counter[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17410_ (.D(_00450_),
    .CLK(clknet_leaf_133_clk),
    .Q(\channels.env_counter[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17411_ (.D(_00451_),
    .CLK(clknet_leaf_134_clk),
    .Q(\channels.env_counter[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17412_ (.D(_00452_),
    .CLK(clknet_leaf_130_clk),
    .Q(\channels.env_counter[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17413_ (.D(_00453_),
    .CLK(clknet_leaf_138_clk),
    .Q(\channels.env_counter[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17414_ (.D(_00454_),
    .CLK(clknet_leaf_139_clk),
    .Q(\channels.env_counter[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17415_ (.D(_00455_),
    .CLK(clknet_leaf_139_clk),
    .Q(\channels.env_counter[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17416_ (.D(_00456_),
    .CLK(clknet_leaf_138_clk),
    .Q(\channels.env_counter[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17417_ (.D(_00457_),
    .CLK(clknet_leaf_153_clk),
    .Q(\channels.env_counter[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17418_ (.D(_00458_),
    .CLK(clknet_leaf_142_clk),
    .Q(\channels.env_counter[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17419_ (.D(_00459_),
    .CLK(clknet_leaf_143_clk),
    .Q(\channels.env_counter[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17420_ (.D(_00460_),
    .CLK(clknet_leaf_151_clk),
    .Q(\channels.env_counter[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17421_ (.D(_00461_),
    .CLK(clknet_leaf_125_clk),
    .Q(\channels.env_counter[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17422_ (.D(_00462_),
    .CLK(clknet_leaf_132_clk),
    .Q(\channels.env_counter[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17423_ (.D(_00463_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.env_counter[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17424_ (.D(_00464_),
    .CLK(clknet_leaf_133_clk),
    .Q(\channels.env_counter[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17425_ (.D(_00465_),
    .CLK(clknet_leaf_134_clk),
    .Q(\channels.env_counter[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17426_ (.D(_00466_),
    .CLK(clknet_leaf_134_clk),
    .Q(\channels.env_counter[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17427_ (.D(_00467_),
    .CLK(clknet_leaf_130_clk),
    .Q(\channels.env_counter[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17428_ (.D(_00468_),
    .CLK(clknet_leaf_136_clk),
    .Q(\channels.env_counter[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17429_ (.D(_00469_),
    .CLK(clknet_leaf_139_clk),
    .Q(\channels.env_counter[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17430_ (.D(_00470_),
    .CLK(clknet_leaf_141_clk),
    .Q(\channels.env_counter[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17431_ (.D(_00471_),
    .CLK(clknet_leaf_140_clk),
    .Q(\channels.env_counter[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17432_ (.D(_00472_),
    .CLK(clknet_leaf_153_clk),
    .Q(\channels.env_counter[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17433_ (.D(_00473_),
    .CLK(clknet_leaf_142_clk),
    .Q(\channels.env_counter[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17434_ (.D(_00474_),
    .CLK(clknet_leaf_142_clk),
    .Q(\channels.env_counter[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17435_ (.D(_00475_),
    .CLK(clknet_leaf_153_clk),
    .Q(\channels.env_counter[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17436_ (.D(_00476_),
    .CLK(clknet_leaf_131_clk),
    .Q(\channels.env_counter[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17437_ (.D(_00477_),
    .CLK(clknet_leaf_125_clk),
    .Q(\channels.env_counter[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17438_ (.D(_00478_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.env_counter[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17439_ (.D(_00479_),
    .CLK(clknet_leaf_171_clk),
    .Q(\channels.adsr_state[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17440_ (.D(_00480_),
    .CLK(clknet_leaf_170_clk),
    .Q(\channels.adsr_state[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17441_ (.D(_00481_),
    .CLK(clknet_leaf_83_clk),
    .Q(\clk_ctr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17442_ (.D(_00482_),
    .CLK(clknet_leaf_80_clk),
    .Q(\clk_ctr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17443_ (.D(_00483_),
    .CLK(clknet_leaf_132_clk),
    .Q(\channels.env_counter[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17444_ (.D(_00484_),
    .CLK(clknet_leaf_135_clk),
    .Q(\channels.env_counter[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17445_ (.D(_00485_),
    .CLK(clknet_leaf_136_clk),
    .Q(\channels.env_counter[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17446_ (.D(_00486_),
    .CLK(clknet_leaf_133_clk),
    .Q(\channels.env_counter[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17447_ (.D(_00487_),
    .CLK(clknet_5_31__leaf_clk),
    .Q(\channels.env_counter[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17448_ (.D(_00488_),
    .CLK(clknet_leaf_140_clk),
    .Q(\channels.env_counter[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17449_ (.D(_00489_),
    .CLK(clknet_leaf_141_clk),
    .Q(\channels.env_counter[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17450_ (.D(_00490_),
    .CLK(clknet_leaf_140_clk),
    .Q(\channels.env_counter[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17451_ (.D(_00491_),
    .CLK(clknet_leaf_153_clk),
    .Q(\channels.env_counter[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17452_ (.D(_00492_),
    .CLK(clknet_leaf_142_clk),
    .Q(\channels.env_counter[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17453_ (.D(_00493_),
    .CLK(clknet_leaf_142_clk),
    .Q(\channels.env_counter[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17454_ (.D(_00494_),
    .CLK(clknet_leaf_152_clk),
    .Q(\channels.env_counter[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17455_ (.D(_00495_),
    .CLK(clknet_leaf_131_clk),
    .Q(\channels.env_counter[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17456_ (.D(_00496_),
    .CLK(clknet_leaf_132_clk),
    .Q(\channels.env_counter[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17457_ (.D(_00497_),
    .CLK(clknet_leaf_130_clk),
    .Q(\channels.env_counter[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17458_ (.D(_00498_),
    .CLK(clknet_leaf_170_clk),
    .Q(\channels.adsr_state[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17459_ (.D(_00499_),
    .CLK(clknet_leaf_170_clk),
    .Q(\channels.adsr_state[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17460_ (.D(_00500_),
    .CLK(clknet_leaf_165_clk),
    .Q(\channels.adsr_state[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17461_ (.D(_00501_),
    .CLK(clknet_leaf_166_clk),
    .Q(\channels.adsr_state[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17462_ (.D(_00502_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.accum[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17463_ (.D(_00503_),
    .CLK(clknet_leaf_184_clk),
    .Q(\channels.accum[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17464_ (.D(_00504_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.accum[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17465_ (.D(_00505_),
    .CLK(clknet_leaf_179_clk),
    .Q(\channels.accum[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17466_ (.D(_00506_),
    .CLK(clknet_leaf_183_clk),
    .Q(\channels.accum[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17467_ (.D(_00507_),
    .CLK(clknet_leaf_173_clk),
    .Q(\channels.accum[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17468_ (.D(_00508_),
    .CLK(clknet_leaf_171_clk),
    .Q(\channels.accum[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17469_ (.D(_00509_),
    .CLK(clknet_leaf_174_clk),
    .Q(\channels.accum[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17470_ (.D(_00510_),
    .CLK(clknet_leaf_150_clk),
    .Q(\channels.accum[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17471_ (.D(_00511_),
    .CLK(clknet_leaf_151_clk),
    .Q(\channels.accum[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17472_ (.D(_00512_),
    .CLK(clknet_leaf_151_clk),
    .Q(\channels.accum[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17473_ (.D(_00513_),
    .CLK(clknet_leaf_149_clk),
    .Q(\channels.accum[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17474_ (.D(_00514_),
    .CLK(clknet_leaf_155_clk),
    .Q(\channels.accum[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17475_ (.D(_00515_),
    .CLK(clknet_leaf_157_clk),
    .Q(\channels.accum[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17476_ (.D(_00516_),
    .CLK(clknet_leaf_159_clk),
    .Q(\channels.accum[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17477_ (.D(_00517_),
    .CLK(clknet_leaf_158_clk),
    .Q(\channels.accum[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17478_ (.D(_00518_),
    .CLK(clknet_leaf_159_clk),
    .Q(\channels.accum[3][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17479_ (.D(_00519_),
    .CLK(clknet_leaf_191_clk),
    .Q(\channels.accum[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17480_ (.D(_00520_),
    .CLK(clknet_leaf_160_clk),
    .Q(\channels.accum[3][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17481_ (.D(_00521_),
    .CLK(clknet_leaf_162_clk),
    .Q(\channels.accum[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17482_ (.D(_00522_),
    .CLK(clknet_leaf_157_clk),
    .Q(\channels.accum[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17483_ (.D(_00523_),
    .CLK(clknet_leaf_194_clk),
    .Q(\channels.accum[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17484_ (.D(_00524_),
    .CLK(clknet_leaf_159_clk),
    .Q(\channels.accum[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17485_ (.D(_00525_),
    .CLK(clknet_leaf_161_clk),
    .Q(\channels.accum[3][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17486_ (.D(_00526_),
    .CLK(clknet_leaf_5_clk),
    .Q(\filters.band[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17487_ (.D(_00527_),
    .CLK(clknet_leaf_4_clk),
    .Q(\filters.band[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17488_ (.D(_00528_),
    .CLK(clknet_leaf_4_clk),
    .Q(\filters.band[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17489_ (.D(_00529_),
    .CLK(clknet_leaf_2_clk),
    .Q(\filters.band[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17490_ (.D(_00530_),
    .CLK(clknet_leaf_0_clk),
    .Q(\filters.band[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17491_ (.D(_00531_),
    .CLK(clknet_leaf_2_clk),
    .Q(\filters.band[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17492_ (.D(_00532_),
    .CLK(clknet_leaf_2_clk),
    .Q(\filters.band[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17493_ (.D(_00533_),
    .CLK(clknet_leaf_2_clk),
    .Q(\filters.band[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17494_ (.D(_00534_),
    .CLK(clknet_leaf_1_clk),
    .Q(\filters.band[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17495_ (.D(_00535_),
    .CLK(clknet_leaf_0_clk),
    .Q(\filters.band[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17496_ (.D(_00536_),
    .CLK(clknet_leaf_245_clk),
    .Q(\filters.band[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17497_ (.D(_00537_),
    .CLK(clknet_leaf_246_clk),
    .Q(\filters.band[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17498_ (.D(_00538_),
    .CLK(clknet_leaf_24_clk),
    .Q(\filters.band[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17499_ (.D(_00539_),
    .CLK(clknet_leaf_246_clk),
    .Q(\filters.band[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17500_ (.D(_00540_),
    .CLK(clknet_leaf_246_clk),
    .Q(\filters.band[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17501_ (.D(_00541_),
    .CLK(clknet_leaf_24_clk),
    .Q(\filters.band[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17502_ (.D(_00542_),
    .CLK(clknet_leaf_27_clk),
    .Q(\filters.band[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17503_ (.D(_00543_),
    .CLK(clknet_leaf_28_clk),
    .Q(\filters.band[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17504_ (.D(_00544_),
    .CLK(clknet_leaf_242_clk),
    .Q(\filters.band[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17505_ (.D(_00545_),
    .CLK(clknet_leaf_242_clk),
    .Q(\filters.band[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17506_ (.D(_00546_),
    .CLK(clknet_leaf_243_clk),
    .Q(\filters.band[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17507_ (.D(_00547_),
    .CLK(clknet_leaf_29_clk),
    .Q(\filters.band[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17508_ (.D(_00548_),
    .CLK(clknet_leaf_29_clk),
    .Q(\filters.band[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17509_ (.D(_00549_),
    .CLK(clknet_leaf_29_clk),
    .Q(\filters.band[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17510_ (.D(_00550_),
    .CLK(clknet_leaf_26_clk),
    .Q(\filters.band[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17511_ (.D(_00551_),
    .CLK(clknet_leaf_30_clk),
    .Q(\filters.band[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17512_ (.D(_00552_),
    .CLK(clknet_leaf_242_clk),
    .Q(\filters.band[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17513_ (.D(_00553_),
    .CLK(clknet_leaf_241_clk),
    .Q(\filters.band[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17514_ (.D(_00554_),
    .CLK(clknet_leaf_241_clk),
    .Q(\filters.band[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17515_ (.D(_00555_),
    .CLK(clknet_leaf_241_clk),
    .Q(\filters.band[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17516_ (.D(_00556_),
    .CLK(clknet_leaf_22_clk),
    .Q(\filters.band[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17517_ (.D(_00557_),
    .CLK(clknet_leaf_26_clk),
    .Q(\filters.band[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17518_ (.D(_00558_),
    .CLK(clknet_leaf_12_clk),
    .Q(\filters.high[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17519_ (.D(_00559_),
    .CLK(clknet_leaf_6_clk),
    .Q(\filters.high[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17520_ (.D(_00560_),
    .CLK(clknet_leaf_6_clk),
    .Q(\filters.high[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17521_ (.D(_00561_),
    .CLK(clknet_leaf_238_clk),
    .Q(\filters.high[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17522_ (.D(_00562_),
    .CLK(clknet_leaf_239_clk),
    .Q(\filters.high[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17523_ (.D(_00563_),
    .CLK(clknet_leaf_7_clk),
    .Q(\filters.high[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17524_ (.D(_00564_),
    .CLK(clknet_leaf_1_clk),
    .Q(\filters.high[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17525_ (.D(_00565_),
    .CLK(clknet_leaf_239_clk),
    .Q(\filters.high[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17526_ (.D(_00566_),
    .CLK(clknet_leaf_238_clk),
    .Q(\filters.high[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17527_ (.D(_00567_),
    .CLK(clknet_leaf_239_clk),
    .Q(\filters.high[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17528_ (.D(_00568_),
    .CLK(clknet_leaf_12_clk),
    .Q(\filters.high[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17529_ (.D(_00569_),
    .CLK(clknet_leaf_11_clk),
    .Q(\filters.high[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17530_ (.D(_00570_),
    .CLK(clknet_leaf_245_clk),
    .Q(\filters.high[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17531_ (.D(_00571_),
    .CLK(clknet_5_6__leaf_clk),
    .Q(\filters.high[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17532_ (.D(_00572_),
    .CLK(clknet_leaf_14_clk),
    .Q(\filters.high[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17533_ (.D(_00573_),
    .CLK(clknet_leaf_23_clk),
    .Q(\filters.high[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17534_ (.D(_00574_),
    .CLK(clknet_leaf_244_clk),
    .Q(\filters.high[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17535_ (.D(_00575_),
    .CLK(clknet_5_1__leaf_clk),
    .Q(\filters.high[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17536_ (.D(_00576_),
    .CLK(clknet_leaf_1_clk),
    .Q(\filters.high[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17537_ (.D(_00577_),
    .CLK(clknet_leaf_244_clk),
    .Q(\filters.high[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17538_ (.D(_00578_),
    .CLK(clknet_leaf_244_clk),
    .Q(\filters.high[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17539_ (.D(_00579_),
    .CLK(clknet_leaf_241_clk),
    .Q(\filters.high[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17540_ (.D(_00580_),
    .CLK(clknet_leaf_245_clk),
    .Q(\filters.high[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17541_ (.D(_00581_),
    .CLK(clknet_leaf_244_clk),
    .Q(\filters.high[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17542_ (.D(_00582_),
    .CLK(clknet_leaf_28_clk),
    .Q(\filters.high[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17543_ (.D(_00583_),
    .CLK(clknet_leaf_23_clk),
    .Q(\filters.high[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17544_ (.D(_00584_),
    .CLK(clknet_leaf_21_clk),
    .Q(\filters.high[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17545_ (.D(_00585_),
    .CLK(clknet_leaf_36_clk),
    .Q(\filters.high[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17546_ (.D(_00586_),
    .CLK(clknet_leaf_22_clk),
    .Q(\filters.high[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17547_ (.D(_00587_),
    .CLK(clknet_leaf_36_clk),
    .Q(\filters.high[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17548_ (.D(_00588_),
    .CLK(clknet_leaf_36_clk),
    .Q(\filters.high[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17549_ (.D(_00589_),
    .CLK(clknet_leaf_21_clk),
    .Q(\filters.high[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17550_ (.D(_00590_),
    .CLK(clknet_leaf_18_clk),
    .Q(\filters.sample_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17551_ (.D(_00591_),
    .CLK(clknet_leaf_18_clk),
    .Q(\filters.sample_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17552_ (.D(_00592_),
    .CLK(clknet_leaf_21_clk),
    .Q(\filters.sample_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17553_ (.D(_00593_),
    .CLK(clknet_leaf_21_clk),
    .Q(\filters.sample_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17554_ (.D(_00594_),
    .CLK(clknet_leaf_21_clk),
    .Q(\filters.sample_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17555_ (.D(_00595_),
    .CLK(clknet_leaf_21_clk),
    .Q(\filters.sample_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17556_ (.D(_00596_),
    .CLK(clknet_leaf_19_clk),
    .Q(\filters.sample_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17557_ (.D(_00597_),
    .CLK(clknet_leaf_19_clk),
    .Q(\filters.sample_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17558_ (.D(_00598_),
    .CLK(clknet_leaf_82_clk),
    .Q(\filters.sample_buff[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17559_ (.D(_00599_),
    .CLK(clknet_leaf_82_clk),
    .Q(\filters.sample_buff[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17560_ (.D(_00600_),
    .CLK(clknet_leaf_82_clk),
    .Q(\filters.sample_buff[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17561_ (.D(_00601_),
    .CLK(clknet_leaf_83_clk),
    .Q(\filters.sample_buff[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17562_ (.D(_00602_),
    .CLK(clknet_leaf_17_clk),
    .Q(\filters.sample_buff[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17563_ (.D(_00603_),
    .CLK(clknet_leaf_85_clk),
    .Q(\filters.sample_buff[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17564_ (.D(_00604_),
    .CLK(clknet_leaf_82_clk),
    .Q(\filters.sample_buff[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17565_ (.D(_00605_),
    .CLK(clknet_leaf_201_clk),
    .Q(\channels.exp_periods[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17566_ (.D(_00606_),
    .CLK(clknet_leaf_201_clk),
    .Q(\channels.exp_periods[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17567_ (.D(_00607_),
    .CLK(clknet_leaf_213_clk),
    .Q(\channels.exp_periods[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17568_ (.D(_00608_),
    .CLK(clknet_leaf_201_clk),
    .Q(\channels.exp_periods[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17569_ (.D(_00609_),
    .CLK(clknet_leaf_201_clk),
    .Q(\channels.exp_periods[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17570_ (.D(_00610_),
    .CLK(clknet_leaf_5_clk),
    .Q(\filters.low[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17571_ (.D(_00611_),
    .CLK(clknet_leaf_5_clk),
    .Q(\filters.low[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17572_ (.D(_00612_),
    .CLK(clknet_leaf_240_clk),
    .Q(\filters.low[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17573_ (.D(_00613_),
    .CLK(clknet_leaf_238_clk),
    .Q(\filters.low[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17574_ (.D(_00614_),
    .CLK(clknet_leaf_0_clk),
    .Q(\filters.low[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17575_ (.D(_00615_),
    .CLK(clknet_leaf_240_clk),
    .Q(\filters.low[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17576_ (.D(_00616_),
    .CLK(clknet_leaf_237_clk),
    .Q(\filters.low[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17577_ (.D(_00617_),
    .CLK(clknet_leaf_179_clk),
    .Q(\filters.low[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17578_ (.D(_00618_),
    .CLK(clknet_leaf_237_clk),
    .Q(\filters.low[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17579_ (.D(_00619_),
    .CLK(clknet_leaf_238_clk),
    .Q(\filters.low[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17580_ (.D(_00620_),
    .CLK(clknet_leaf_6_clk),
    .Q(\filters.low[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17581_ (.D(_00621_),
    .CLK(clknet_leaf_13_clk),
    .Q(\filters.low[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17582_ (.D(_00622_),
    .CLK(clknet_leaf_13_clk),
    .Q(\filters.low[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17583_ (.D(_00623_),
    .CLK(clknet_leaf_23_clk),
    .Q(\filters.low[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17584_ (.D(_00624_),
    .CLK(clknet_leaf_23_clk),
    .Q(\filters.low[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17585_ (.D(_00625_),
    .CLK(clknet_leaf_24_clk),
    .Q(\filters.low[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17586_ (.D(_00626_),
    .CLK(clknet_leaf_26_clk),
    .Q(\filters.low[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17587_ (.D(_00627_),
    .CLK(clknet_leaf_28_clk),
    .Q(\filters.low[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17588_ (.D(_00628_),
    .CLK(clknet_leaf_242_clk),
    .Q(\filters.low[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17589_ (.D(_00629_),
    .CLK(clknet_leaf_242_clk),
    .Q(\filters.low[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17590_ (.D(_00630_),
    .CLK(clknet_leaf_242_clk),
    .Q(\filters.low[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17591_ (.D(_00631_),
    .CLK(clknet_leaf_243_clk),
    .Q(\filters.low[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17592_ (.D(_00632_),
    .CLK(clknet_leaf_30_clk),
    .Q(\filters.low[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17593_ (.D(_00633_),
    .CLK(clknet_5_2__leaf_clk),
    .Q(\filters.low[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17594_ (.D(_00634_),
    .CLK(clknet_leaf_27_clk),
    .Q(\filters.low[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17595_ (.D(_00635_),
    .CLK(clknet_leaf_33_clk),
    .Q(\filters.low[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17596_ (.D(_00636_),
    .CLK(clknet_leaf_33_clk),
    .Q(\filters.low[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17597_ (.D(_00637_),
    .CLK(clknet_leaf_33_clk),
    .Q(\filters.low[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17598_ (.D(_00638_),
    .CLK(clknet_5_2__leaf_clk),
    .Q(\filters.low[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17599_ (.D(_00639_),
    .CLK(clknet_leaf_33_clk),
    .Q(\filters.low[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17600_ (.D(_00640_),
    .CLK(clknet_leaf_22_clk),
    .Q(\filters.low[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17601_ (.D(_00641_),
    .CLK(clknet_leaf_26_clk),
    .Q(\filters.low[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17602_ (.D(_00642_),
    .CLK(clknet_5_4__leaf_clk),
    .Q(\filters.filter_step[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _17603_ (.D(_00643_),
    .CLK(clknet_leaf_3_clk),
    .Q(\filters.filter_step[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17604_ (.D(_00644_),
    .CLK(clknet_leaf_3_clk),
    .Q(\filters.filter_step[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17605_ (.D(_00645_),
    .CLK(clknet_leaf_37_clk),
    .Q(\spi_dac_i.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17606_ (.D(_00646_),
    .CLK(clknet_leaf_36_clk),
    .Q(\spi_dac_i.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17607_ (.D(_00647_),
    .CLK(clknet_leaf_36_clk),
    .Q(\spi_dac_i.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17608_ (.D(_00648_),
    .CLK(clknet_leaf_36_clk),
    .Q(\spi_dac_i.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17609_ (.D(_00649_),
    .CLK(clknet_leaf_21_clk),
    .Q(\spi_dac_i.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17610_ (.D(_00650_),
    .CLK(clknet_leaf_36_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17611_ (.D(_00651_),
    .CLK(clknet_leaf_34_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17612_ (.D(_00652_),
    .CLK(clknet_leaf_34_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17613_ (.D(_00653_),
    .CLK(clknet_leaf_34_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17614_ (.D(_00654_),
    .CLK(clknet_leaf_34_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17615_ (.D(_00655_),
    .CLK(clknet_leaf_34_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17616_ (.D(_00656_),
    .CLK(clknet_leaf_35_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17617_ (.D(_00657_),
    .CLK(clknet_leaf_35_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17618_ (.D(_00658_),
    .CLK(clknet_leaf_35_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17619_ (.D(_00659_),
    .CLK(clknet_leaf_39_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17620_ (.D(_00660_),
    .CLK(clknet_leaf_39_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17621_ (.D(_00661_),
    .CLK(clknet_leaf_38_clk),
    .Q(\spi_dac_i.spi_dat_buff_1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17622_ (.D(_00662_),
    .CLK(clknet_leaf_37_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17623_ (.D(_00663_),
    .CLK(clknet_leaf_37_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17624_ (.D(_00664_),
    .CLK(clknet_leaf_20_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17625_ (.D(_00665_),
    .CLK(clknet_leaf_20_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17626_ (.D(_00666_),
    .CLK(clknet_leaf_19_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17627_ (.D(_00667_),
    .CLK(clknet_leaf_82_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17628_ (.D(_00668_),
    .CLK(clknet_leaf_81_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17629_ (.D(_00669_),
    .CLK(clknet_leaf_81_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17630_ (.D(_00670_),
    .CLK(clknet_leaf_56_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17631_ (.D(_00671_),
    .CLK(clknet_leaf_56_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17632_ (.D(_00672_),
    .CLK(clknet_leaf_38_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17633_ (.D(_00673_),
    .CLK(clknet_leaf_38_clk),
    .Q(\spi_dac_i.spi_dat_buff_0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17634_ (.D(_00674_),
    .CLK(clknet_leaf_38_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17635_ (.D(_00675_),
    .CLK(clknet_leaf_38_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17636_ (.D(_00676_),
    .CLK(clknet_leaf_44_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17637_ (.D(_00677_),
    .CLK(clknet_leaf_166_clk),
    .Q(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17638_ (.D(_00678_),
    .CLK(clknet_leaf_169_clk),
    .Q(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17639_ (.D(_00679_),
    .CLK(clknet_leaf_133_clk),
    .Q(\channels.env_counter[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17640_ (.D(_00680_),
    .CLK(clknet_leaf_135_clk),
    .Q(\channels.env_counter[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17641_ (.D(_00681_),
    .CLK(clknet_leaf_135_clk),
    .Q(\channels.env_counter[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17642_ (.D(_00682_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.env_counter[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17643_ (.D(_00683_),
    .CLK(clknet_leaf_138_clk),
    .Q(\channels.env_counter[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17644_ (.D(_00684_),
    .CLK(clknet_leaf_141_clk),
    .Q(\channels.env_counter[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17645_ (.D(_00685_),
    .CLK(clknet_leaf_141_clk),
    .Q(\channels.env_counter[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17646_ (.D(_00686_),
    .CLK(clknet_leaf_136_clk),
    .Q(\channels.env_counter[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17647_ (.D(_00687_),
    .CLK(clknet_leaf_154_clk),
    .Q(\channels.env_counter[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17648_ (.D(_00688_),
    .CLK(clknet_leaf_141_clk),
    .Q(\channels.env_counter[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17649_ (.D(_00689_),
    .CLK(clknet_leaf_145_clk),
    .Q(\channels.env_counter[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17650_ (.D(_00690_),
    .CLK(clknet_leaf_151_clk),
    .Q(\channels.env_counter[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17651_ (.D(_00691_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.env_counter[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17652_ (.D(_00692_),
    .CLK(clknet_leaf_136_clk),
    .Q(\channels.env_counter[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17653_ (.D(_00693_),
    .CLK(clknet_leaf_129_clk),
    .Q(\channels.env_counter[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17654_ (.D(_00694_),
    .CLK(clknet_leaf_185_clk),
    .Q(\channels.env_vol[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17655_ (.D(_00695_),
    .CLK(clknet_leaf_208_clk),
    .Q(\channels.env_vol[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17656_ (.D(_00696_),
    .CLK(clknet_leaf_207_clk),
    .Q(\channels.env_vol[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17657_ (.D(_00697_),
    .CLK(clknet_leaf_207_clk),
    .Q(\channels.env_vol[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17658_ (.D(_00698_),
    .CLK(clknet_leaf_212_clk),
    .Q(\channels.env_vol[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17659_ (.D(_00699_),
    .CLK(clknet_leaf_207_clk),
    .Q(\channels.env_vol[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17660_ (.D(_00700_),
    .CLK(clknet_leaf_212_clk),
    .Q(\channels.env_vol[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17661_ (.D(_00701_),
    .CLK(clknet_leaf_204_clk),
    .Q(\channels.env_vol[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17662_ (.D(_00702_),
    .CLK(clknet_leaf_195_clk),
    .Q(\channels.exp_counter[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17663_ (.D(_00703_),
    .CLK(clknet_leaf_195_clk),
    .Q(\channels.exp_counter[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17664_ (.D(_00704_),
    .CLK(clknet_leaf_197_clk),
    .Q(\channels.exp_counter[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17665_ (.D(_00705_),
    .CLK(clknet_leaf_199_clk),
    .Q(\channels.exp_counter[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17666_ (.D(_00706_),
    .CLK(clknet_leaf_192_clk),
    .Q(\channels.exp_counter[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17667_ (.D(_00707_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.ch3_env[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17668_ (.D(_00708_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.ch3_env[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17669_ (.D(_00709_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.ch3_env[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17670_ (.D(_00710_),
    .CLK(clknet_leaf_186_clk),
    .Q(\channels.ch3_env[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17671_ (.D(_00711_),
    .CLK(clknet_leaf_204_clk),
    .Q(\channels.ch3_env[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17672_ (.D(_00712_),
    .CLK(clknet_leaf_205_clk),
    .Q(\channels.ch3_env[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17673_ (.D(_00713_),
    .CLK(clknet_5_22__leaf_clk),
    .Q(\channels.ch3_env[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17674_ (.D(_00714_),
    .CLK(clknet_leaf_199_clk),
    .Q(\channels.ch3_env[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17675_ (.D(_00715_),
    .CLK(clknet_leaf_43_clk),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17676_ (.D(_00716_),
    .CLK(clknet_leaf_43_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17677_ (.D(_00717_),
    .CLK(clknet_leaf_43_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17678_ (.D(_00718_),
    .CLK(clknet_leaf_43_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17679_ (.D(_00719_),
    .CLK(clknet_leaf_43_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17680_ (.D(_00720_),
    .CLK(clknet_leaf_44_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17681_ (.D(_00721_),
    .CLK(clknet_leaf_44_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17682_ (.D(_00722_),
    .CLK(clknet_leaf_44_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17683_ (.D(_00723_),
    .CLK(clknet_leaf_45_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17684_ (.D(_00724_),
    .CLK(clknet_leaf_45_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17685_ (.D(_00725_),
    .CLK(clknet_leaf_47_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17686_ (.D(_00726_),
    .CLK(clknet_leaf_47_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17687_ (.D(_00727_),
    .CLK(clknet_leaf_45_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17688_ (.D(_00728_),
    .CLK(clknet_leaf_45_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17689_ (.D(_00729_),
    .CLK(clknet_leaf_43_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.lfsr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17690_ (.D(_00730_),
    .CLK(clknet_leaf_55_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17691_ (.D(_00731_),
    .CLK(clknet_leaf_56_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17692_ (.D(_00732_),
    .CLK(clknet_leaf_55_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17693_ (.D(_00733_),
    .CLK(clknet_leaf_55_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17694_ (.D(_00734_),
    .CLK(clknet_leaf_54_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17695_ (.D(_00735_),
    .CLK(clknet_leaf_52_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17696_ (.D(_00736_),
    .CLK(clknet_leaf_55_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17697_ (.D(_00737_),
    .CLK(clknet_leaf_47_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17698_ (.D(_00738_),
    .CLK(clknet_leaf_61_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17699_ (.D(_00739_),
    .CLK(clknet_leaf_49_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17700_ (.D(_00740_),
    .CLK(clknet_leaf_47_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17701_ (.D(_00741_),
    .CLK(clknet_leaf_47_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17702_ (.D(_00742_),
    .CLK(clknet_leaf_47_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17703_ (.D(_00743_),
    .CLK(clknet_leaf_48_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17704_ (.D(_00744_),
    .CLK(clknet_leaf_48_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17705_ (.D(_00745_),
    .CLK(clknet_leaf_50_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17706_ (.D(_00746_),
    .CLK(clknet_leaf_49_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17707_ (.D(_00747_),
    .CLK(clknet_leaf_50_clk),
    .Q(\tt_um_rejunity_sn76489.tone[2].gen.counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17708_ (.D(_00748_),
    .CLK(clknet_leaf_53_clk),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17709_ (.D(_00749_),
    .CLK(clknet_leaf_62_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17710_ (.D(_00750_),
    .CLK(clknet_leaf_62_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17711_ (.D(_00751_),
    .CLK(clknet_leaf_62_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17712_ (.D(_00752_),
    .CLK(clknet_leaf_63_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17713_ (.D(_00753_),
    .CLK(clknet_leaf_61_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17714_ (.D(_00754_),
    .CLK(clknet_leaf_61_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17715_ (.D(_00755_),
    .CLK(clknet_leaf_61_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17716_ (.D(_00756_),
    .CLK(clknet_leaf_64_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17717_ (.D(_00757_),
    .CLK(clknet_leaf_60_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17718_ (.D(_00758_),
    .CLK(clknet_leaf_60_clk),
    .Q(\tt_um_rejunity_sn76489.tone[1].gen.counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17719_ (.D(_00759_),
    .CLK(clknet_leaf_51_clk),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17720_ (.D(_00760_),
    .CLK(clknet_leaf_214_clk),
    .Q(\channels.lfsr[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17721_ (.D(_00761_),
    .CLK(clknet_leaf_215_clk),
    .Q(\channels.lfsr[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17722_ (.D(_00762_),
    .CLK(clknet_leaf_216_clk),
    .Q(\channels.lfsr[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17723_ (.D(_00763_),
    .CLK(clknet_leaf_216_clk),
    .Q(\channels.lfsr[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17724_ (.D(_00764_),
    .CLK(clknet_leaf_218_clk),
    .Q(\channels.lfsr[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17725_ (.D(_00765_),
    .CLK(clknet_leaf_218_clk),
    .Q(\channels.lfsr[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17726_ (.D(_00766_),
    .CLK(clknet_leaf_220_clk),
    .Q(\channels.lfsr[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17727_ (.D(_00767_),
    .CLK(clknet_leaf_220_clk),
    .Q(\channels.lfsr[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17728_ (.D(_00768_),
    .CLK(clknet_leaf_221_clk),
    .Q(\channels.lfsr[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17729_ (.D(_00769_),
    .CLK(clknet_leaf_223_clk),
    .Q(\channels.lfsr[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17730_ (.D(_00770_),
    .CLK(clknet_leaf_222_clk),
    .Q(\channels.lfsr[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17731_ (.D(_00771_),
    .CLK(clknet_leaf_225_clk),
    .Q(\channels.lfsr[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17732_ (.D(_00772_),
    .CLK(clknet_leaf_227_clk),
    .Q(\channels.lfsr[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17733_ (.D(_00773_),
    .CLK(clknet_leaf_228_clk),
    .Q(\channels.lfsr[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17734_ (.D(_00774_),
    .CLK(clknet_leaf_228_clk),
    .Q(\channels.lfsr[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17735_ (.D(_00775_),
    .CLK(clknet_leaf_234_clk),
    .Q(\channels.lfsr[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17736_ (.D(_00776_),
    .CLK(clknet_leaf_233_clk),
    .Q(\channels.lfsr[0][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17737_ (.D(_00777_),
    .CLK(clknet_leaf_229_clk),
    .Q(\channels.lfsr[0][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17738_ (.D(_00778_),
    .CLK(clknet_leaf_229_clk),
    .Q(\channels.lfsr[0][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17739_ (.D(_00779_),
    .CLK(clknet_leaf_232_clk),
    .Q(\channels.lfsr[0][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17740_ (.D(_00780_),
    .CLK(clknet_leaf_231_clk),
    .Q(\channels.lfsr[0][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17741_ (.D(_00781_),
    .CLK(clknet_leaf_224_clk),
    .Q(\channels.lfsr[0][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17742_ (.D(_00782_),
    .CLK(clknet_leaf_224_clk),
    .Q(\channels.lfsr[0][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17743_ (.D(_00783_),
    .CLK(clknet_leaf_64_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17744_ (.D(_00784_),
    .CLK(clknet_leaf_63_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17745_ (.D(_00785_),
    .CLK(clknet_leaf_66_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17746_ (.D(_00786_),
    .CLK(clknet_leaf_66_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17747_ (.D(_00787_),
    .CLK(clknet_leaf_65_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17748_ (.D(_00788_),
    .CLK(clknet_leaf_71_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17749_ (.D(_00789_),
    .CLK(clknet_leaf_71_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17750_ (.D(_00790_),
    .CLK(clknet_leaf_65_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17751_ (.D(_00791_),
    .CLK(clknet_leaf_64_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17752_ (.D(_00792_),
    .CLK(clknet_leaf_59_clk),
    .Q(\tt_um_rejunity_sn76489.tone[0].gen.counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17753_ (.D(_00793_),
    .CLK(clknet_leaf_50_clk),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.in ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17754_ (.D(_00794_),
    .CLK(clknet_leaf_53_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17755_ (.D(_00795_),
    .CLK(clknet_leaf_53_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17756_ (.D(_00796_),
    .CLK(clknet_leaf_50_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17757_ (.D(_00797_),
    .CLK(clknet_leaf_50_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17758_ (.D(_00798_),
    .CLK(clknet_leaf_58_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17759_ (.D(_00799_),
    .CLK(clknet_leaf_54_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17760_ (.D(_00800_),
    .CLK(clknet_leaf_58_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17761_ (.D(_00801_),
    .CLK(clknet_leaf_58_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17762_ (.D(_00802_),
    .CLK(clknet_leaf_60_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17763_ (.D(_00803_),
    .CLK(clknet_leaf_60_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17764_ (.D(_00804_),
    .CLK(clknet_leaf_58_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17765_ (.D(_00805_),
    .CLK(clknet_leaf_60_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17766_ (.D(_00806_),
    .CLK(clknet_leaf_72_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17767_ (.D(_00807_),
    .CLK(clknet_5_14__leaf_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17768_ (.D(_00808_),
    .CLK(clknet_leaf_59_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17769_ (.D(_00809_),
    .CLK(clknet_leaf_59_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17770_ (.D(_00810_),
    .CLK(clknet_leaf_59_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17771_ (.D(_00811_),
    .CLK(clknet_leaf_59_clk),
    .Q(\tt_um_rejunity_sn76489.control_tone_freq[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17772_ (.D(_00812_),
    .CLK(clknet_leaf_41_clk),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17773_ (.D(_00813_),
    .CLK(clknet_leaf_41_clk),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17774_ (.D(_00814_),
    .CLK(clknet_leaf_41_clk),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17775_ (.D(_00815_),
    .CLK(clknet_5_8__leaf_clk),
    .Q(\tt_um_rejunity_sn76489.chan[3].attenuation.control[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17776_ (.D(_00816_),
    .CLK(clknet_leaf_52_clk),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17777_ (.D(_00817_),
    .CLK(clknet_leaf_40_clk),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _17778_ (.D(_00818_),
    .CLK(clknet_leaf_40_clk),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17779_ (.D(_00819_),
    .CLK(clknet_leaf_40_clk),
    .Q(\tt_um_rejunity_sn76489.chan[2].attenuation.control[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17780_ (.D(_00820_),
    .CLK(clknet_leaf_46_clk),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17781_ (.D(_00821_),
    .CLK(clknet_leaf_46_clk),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17782_ (.D(_00822_),
    .CLK(clknet_leaf_46_clk),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17783_ (.D(_00823_),
    .CLK(clknet_leaf_46_clk),
    .Q(\tt_um_rejunity_sn76489.chan[1].attenuation.control[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17784_ (.D(_00824_),
    .CLK(clknet_leaf_52_clk),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17785_ (.D(_00825_),
    .CLK(clknet_leaf_51_clk),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17786_ (.D(_00826_),
    .CLK(clknet_leaf_51_clk),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17787_ (.D(_00827_),
    .CLK(clknet_leaf_51_clk),
    .Q(\tt_um_rejunity_sn76489.chan[0].attenuation.control[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17788_ (.D(_00828_),
    .CLK(clknet_leaf_57_clk),
    .Q(\tt_um_rejunity_sn76489.noise[0].gen.restart_noise ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17789_ (.D(_00829_),
    .CLK(clknet_leaf_80_clk),
    .Q(\tt_um_rejunity_sn76489.latch_control_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17790_ (.D(_00830_),
    .CLK(clknet_leaf_80_clk),
    .Q(\tt_um_rejunity_sn76489.latch_control_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17791_ (.D(_00831_),
    .CLK(clknet_leaf_80_clk),
    .Q(\tt_um_rejunity_sn76489.latch_control_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17792_ (.D(_00832_),
    .CLK(clknet_leaf_80_clk),
    .Q(\tt_um_rejunity_sn76489.clk_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17793_ (.D(_00833_),
    .CLK(clknet_leaf_81_clk),
    .Q(\tt_um_rejunity_sn76489.clk_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17794_ (.D(_00834_),
    .CLK(clknet_leaf_81_clk),
    .Q(\tt_um_rejunity_sn76489.clk_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17795_ (.D(_00835_),
    .CLK(clknet_leaf_81_clk),
    .Q(\tt_um_rejunity_sn76489.clk_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17796_ (.D(_00836_),
    .CLK(clknet_leaf_57_clk),
    .Q(\tt_um_rejunity_sn76489.clk_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17797_ (.D(_00837_),
    .CLK(clknet_leaf_200_clk),
    .Q(\channels.exp_periods[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17798_ (.D(_00838_),
    .CLK(clknet_leaf_202_clk),
    .Q(\channels.exp_periods[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17799_ (.D(_00839_),
    .CLK(clknet_leaf_212_clk),
    .Q(\channels.exp_periods[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17800_ (.D(_00840_),
    .CLK(clknet_leaf_203_clk),
    .Q(\channels.exp_periods[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17801_ (.D(_00841_),
    .CLK(clknet_leaf_205_clk),
    .Q(\channels.exp_periods[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17802_ (.D(_00842_),
    .CLK(clknet_leaf_200_clk),
    .Q(\channels.exp_periods[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17803_ (.D(_00843_),
    .CLK(clknet_leaf_203_clk),
    .Q(\channels.exp_periods[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17804_ (.D(_00844_),
    .CLK(clknet_leaf_202_clk),
    .Q(\channels.exp_periods[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17805_ (.D(_00845_),
    .CLK(clknet_leaf_205_clk),
    .Q(\channels.exp_periods[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17806_ (.D(_00846_),
    .CLK(clknet_leaf_199_clk),
    .Q(\channels.exp_periods[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17807_ (.D(_00847_),
    .CLK(clknet_leaf_195_clk),
    .Q(\channels.exp_counter[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17808_ (.D(_00848_),
    .CLK(clknet_leaf_195_clk),
    .Q(\channels.exp_counter[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17809_ (.D(_00849_),
    .CLK(clknet_leaf_197_clk),
    .Q(\channels.exp_counter[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17810_ (.D(_00850_),
    .CLK(clknet_leaf_197_clk),
    .Q(\channels.exp_counter[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17811_ (.D(_00851_),
    .CLK(clknet_leaf_191_clk),
    .Q(\channels.exp_counter[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17812_ (.D(_00852_),
    .CLK(clknet_leaf_200_clk),
    .Q(\channels.exp_periods[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17813_ (.D(_00853_),
    .CLK(clknet_leaf_212_clk),
    .Q(\channels.exp_periods[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17814_ (.D(_00854_),
    .CLK(clknet_leaf_213_clk),
    .Q(\channels.exp_periods[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17815_ (.D(_00855_),
    .CLK(clknet_leaf_204_clk),
    .Q(\channels.exp_periods[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17816_ (.D(_00856_),
    .CLK(clknet_leaf_205_clk),
    .Q(\channels.exp_periods[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17817_ (.D(_00857_),
    .CLK(clknet_leaf_54_clk),
    .Q(\tt_um_rejunity_sn76489.control_noise[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17818_ (.D(_00858_),
    .CLK(clknet_leaf_57_clk),
    .Q(\tt_um_rejunity_sn76489.control_noise[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _17819_ (.D(_00859_),
    .CLK(clknet_leaf_53_clk),
    .Q(\tt_um_rejunity_sn76489.control_noise[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_3_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_0__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_10__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_10__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_11__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_11__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_12__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_12__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_13__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_13__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_14__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_14__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_15__f_clk (.I(clknet_3_3_0_clk),
    .Z(clknet_5_15__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_16__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_16__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_17__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_17__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_18__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_18__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_19__f_clk (.I(clknet_3_4_0_clk),
    .Z(clknet_5_19__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_1__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_20__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_20__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_21__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_21__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_22__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_22__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_23__f_clk (.I(clknet_3_5_0_clk),
    .Z(clknet_5_23__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_24__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_24__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_25__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_25__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_26__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_26__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_27__f_clk (.I(clknet_3_6_0_clk),
    .Z(clknet_5_27__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_28__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_28__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_29__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_29__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_2__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_30__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_30__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_31__f_clk (.I(clknet_3_7_0_clk),
    .Z(clknet_5_31__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_3__f_clk (.I(clknet_3_0_0_clk),
    .Z(clknet_5_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_4__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_4__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_5__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_5__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_6__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_6__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_7__f_clk (.I(clknet_3_1_0_clk),
    .Z(clknet_5_7__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_8__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_8__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_5_9__f_clk (.I(clknet_3_2_0_clk),
    .Z(clknet_5_9__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_111_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_116_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_117_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_118_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_119_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_120_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_clk (.I(clknet_5_26__leaf_clk),
    .Z(clknet_leaf_121_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_123_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_124_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_125_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_126_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_127_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_128_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_129_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_130_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_131_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_131_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_132_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_133_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_133_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_134_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_135_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_136_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_136_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_138_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_138_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_139_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_139_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_140_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_140_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_141_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_141_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_142_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_142_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_143_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_143_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_144_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_144_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_145_clk (.I(clknet_5_30__leaf_clk),
    .Z(clknet_leaf_145_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_146_clk (.I(clknet_5_27__leaf_clk),
    .Z(clknet_leaf_146_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_147_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_147_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_148_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_148_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_149_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_149_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_150_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_150_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_151_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_151_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_152_clk (.I(clknet_5_31__leaf_clk),
    .Z(clknet_leaf_152_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_153_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_153_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_154_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_154_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_155_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_155_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_156_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_156_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_157_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_157_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_158_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_158_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_159_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_159_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_160_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_160_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_161_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_161_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_162_clk (.I(clknet_5_29__leaf_clk),
    .Z(clknet_leaf_162_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_163_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_163_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_164_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_164_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_165_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_165_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_166_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_166_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_167_clk (.I(clknet_5_28__leaf_clk),
    .Z(clknet_leaf_167_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_168_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_168_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_169_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_169_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_170_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_170_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_171_clk (.I(clknet_5_25__leaf_clk),
    .Z(clknet_leaf_171_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_172_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_172_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_173_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_173_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_174_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_174_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_175_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_175_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_176_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_176_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_177_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_177_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_178_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_178_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_179_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_179_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_180_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_180_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_181_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_181_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_183_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_183_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_184_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_184_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_185_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_185_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_186_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_186_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_187_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_187_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_188_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_188_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_190_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_190_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_191_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_191_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_192_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_192_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_193_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_193_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_194_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_194_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_195_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_195_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_196_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_196_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_197_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_197_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_199_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_199_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clk (.I(clknet_5_6__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_200_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_200_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_201_clk (.I(clknet_5_23__leaf_clk),
    .Z(clknet_leaf_201_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_202_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_202_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_203_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_203_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_204_clk (.I(clknet_5_22__leaf_clk),
    .Z(clknet_leaf_204_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_205_clk (.I(clknet_5_19__leaf_clk),
    .Z(clknet_leaf_205_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_207_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_207_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_208_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_208_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_209_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_209_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_210_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_210_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_211_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_211_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_212_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_212_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_213_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_213_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_214_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_214_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_215_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_215_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_216_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_216_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_217_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_217_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_218_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_218_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_219_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_219_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_220_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_220_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_221_clk (.I(clknet_5_21__leaf_clk),
    .Z(clknet_leaf_221_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_222_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_222_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_223_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_223_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_224_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_224_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_225_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_225_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_226_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_226_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_227_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_227_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_228_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_228_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_229_clk (.I(clknet_5_17__leaf_clk),
    .Z(clknet_leaf_229_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_230_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_230_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_231_clk (.I(clknet_5_20__leaf_clk),
    .Z(clknet_leaf_231_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_232_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_232_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_233_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_233_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_234_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_234_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_235_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_235_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_236_clk (.I(clknet_5_16__leaf_clk),
    .Z(clknet_leaf_236_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_237_clk (.I(clknet_5_18__leaf_clk),
    .Z(clknet_leaf_237_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_238_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_238_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_239_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_239_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_240_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_240_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_241_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_241_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_242_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_242_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_243_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_243_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_244_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_244_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_245_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_245_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_246_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_246_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clk (.I(clknet_5_0__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_5_1__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clk (.I(clknet_5_2__leaf_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clk (.I(clknet_5_3__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_clk (.I(clknet_5_10__leaf_clk),
    .Z(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clk (.I(clknet_5_8__leaf_clk),
    .Z(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_clk (.I(clknet_5_11__leaf_clk),
    .Z(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_5_4__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_clk (.I(clknet_5_14__leaf_clk),
    .Z(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_clk (.I(clknet_5_15__leaf_clk),
    .Z(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_clk (.I(clknet_5_9__leaf_clk),
    .Z(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_clk (.I(clknet_5_12__leaf_clk),
    .Z(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_89_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_95_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_clk (.I(clknet_5_7__leaf_clk),
    .Z(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_clk (.I(clknet_5_24__leaf_clk),
    .Z(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_clk (.I(clknet_5_13__leaf_clk),
    .Z(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clk (.I(clknet_5_5__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1 (.I(addr[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input10 (.I(bus_in[3]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(bus_in[4]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input12 (.I(bus_in[5]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input13 (.I(bus_in[6]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input14 (.I(bus_in[7]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(bus_we),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input16 (.I(rst),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input2 (.I(addr[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(addr[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input4 (.I(addr[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input5 (.I(addr[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(bus_cyc),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input7 (.I(bus_in[0]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input8 (.I(bus_in[1]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input9 (.I(bus_in[2]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output17 (.I(net17),
    .Z(DAC_clk));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output18 (.I(net18),
    .Z(DAC_dat_1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output19 (.I(net19),
    .Z(DAC_dat_2));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(DAC_le));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(bus_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(bus_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(bus_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(bus_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output25 (.I(net25),
    .Z(bus_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output26 (.I(net26),
    .Z(bus_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output27 (.I(net27),
    .Z(bus_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output28 (.I(net28),
    .Z(bus_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 rebuffer1 (.I(_07380_),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer10 (.I(_05057_),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer11 (.I(_05404_),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer12 (.I(_05313_),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer13 (.I(_05180_),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer14 (.I(_05452_),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer15 (.I(_04415_),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer16 (.I(net43),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer17 (.I(_05373_),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer18 (.I(_05196_),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer19 (.I(_04388_),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer2 (.I(_06536_),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer20 (.I(_04268_),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer21 (.I(net48),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer22 (.I(net51),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer23 (.I(net71),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer24 (.I(_05221_),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer25 (.I(_04301_),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer26 (.I(_03399_),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer27 (.I(net54),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer28 (.I(_04246_),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 rebuffer29 (.I(_04897_),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 rebuffer3 (.I(_06859_),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer30 (.I(_04190_),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer31 (.I(_04205_),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer32 (.I(_04416_),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer33 (.I(_05357_),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer34 (.I(_05429_),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer35 (.I(_04257_),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer36 (.I(_05255_),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer37 (.I(_05063_),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer38 (.I(_04843_),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer39 (.I(_04519_),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer4 (.I(_06628_),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer40 (.I(_04222_),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer41 (.I(_03288_),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer42 (.I(_04205_),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlya_1 rebuffer43 (.I(_07380_),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(_04194_),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer6 (.I(_04194_),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer7 (.I(net42),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer8 (.I(_05460_),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer9 (.I(_04377_),
    .Z(net37));
endmodule

