magic
tech gf180mcuD
magscale 1 5
timestamp 1701123629
<< obsm1 >>
rect 672 1538 104328 68238
<< metal2 >>
rect 672 69600 728 70000
rect 2016 69600 2072 70000
rect 3360 69600 3416 70000
rect 4704 69600 4760 70000
rect 6048 69600 6104 70000
rect 7392 69600 7448 70000
rect 8736 69600 8792 70000
rect 10080 69600 10136 70000
rect 11424 69600 11480 70000
rect 12768 69600 12824 70000
rect 14112 69600 14168 70000
rect 15456 69600 15512 70000
rect 16800 69600 16856 70000
rect 18144 69600 18200 70000
rect 19488 69600 19544 70000
rect 20832 69600 20888 70000
rect 22176 69600 22232 70000
rect 23520 69600 23576 70000
rect 24864 69600 24920 70000
rect 26208 69600 26264 70000
rect 27552 69600 27608 70000
rect 28896 69600 28952 70000
rect 30240 69600 30296 70000
rect 31584 69600 31640 70000
rect 32928 69600 32984 70000
rect 34272 69600 34328 70000
rect 35616 69600 35672 70000
rect 36960 69600 37016 70000
rect 38304 69600 38360 70000
rect 39648 69600 39704 70000
rect 40992 69600 41048 70000
rect 42336 69600 42392 70000
rect 43680 69600 43736 70000
rect 45024 69600 45080 70000
rect 46368 69600 46424 70000
rect 47712 69600 47768 70000
rect 49056 69600 49112 70000
rect 50400 69600 50456 70000
rect 51744 69600 51800 70000
rect 53088 69600 53144 70000
rect 54432 69600 54488 70000
rect 55776 69600 55832 70000
rect 57120 69600 57176 70000
rect 58464 69600 58520 70000
rect 59808 69600 59864 70000
rect 61152 69600 61208 70000
rect 62496 69600 62552 70000
rect 63840 69600 63896 70000
rect 65184 69600 65240 70000
rect 66528 69600 66584 70000
rect 67872 69600 67928 70000
rect 69216 69600 69272 70000
rect 70560 69600 70616 70000
rect 71904 69600 71960 70000
rect 73248 69600 73304 70000
rect 74592 69600 74648 70000
rect 75936 69600 75992 70000
rect 77280 69600 77336 70000
rect 78624 69600 78680 70000
rect 79968 69600 80024 70000
rect 81312 69600 81368 70000
rect 82656 69600 82712 70000
rect 84000 69600 84056 70000
rect 85344 69600 85400 70000
rect 86688 69600 86744 70000
rect 88032 69600 88088 70000
rect 89376 69600 89432 70000
rect 90720 69600 90776 70000
rect 92064 69600 92120 70000
rect 93408 69600 93464 70000
rect 94752 69600 94808 70000
rect 96096 69600 96152 70000
rect 97440 69600 97496 70000
rect 98784 69600 98840 70000
rect 100128 69600 100184 70000
rect 101472 69600 101528 70000
rect 102816 69600 102872 70000
rect 104160 69600 104216 70000
rect 1568 0 1624 400
rect 2576 0 2632 400
rect 3584 0 3640 400
rect 4592 0 4648 400
rect 5600 0 5656 400
rect 6608 0 6664 400
rect 7616 0 7672 400
rect 8624 0 8680 400
rect 9632 0 9688 400
rect 10640 0 10696 400
rect 11648 0 11704 400
rect 12656 0 12712 400
rect 13664 0 13720 400
rect 14672 0 14728 400
rect 15680 0 15736 400
rect 16688 0 16744 400
rect 17696 0 17752 400
rect 18704 0 18760 400
rect 19712 0 19768 400
rect 20720 0 20776 400
rect 21728 0 21784 400
rect 22736 0 22792 400
rect 23744 0 23800 400
rect 24752 0 24808 400
rect 25760 0 25816 400
rect 26768 0 26824 400
rect 27776 0 27832 400
rect 28784 0 28840 400
rect 29792 0 29848 400
rect 30800 0 30856 400
rect 31808 0 31864 400
rect 32816 0 32872 400
rect 33824 0 33880 400
rect 34832 0 34888 400
rect 35840 0 35896 400
rect 36848 0 36904 400
rect 37856 0 37912 400
rect 38864 0 38920 400
rect 39872 0 39928 400
rect 40880 0 40936 400
rect 41888 0 41944 400
rect 42896 0 42952 400
rect 43904 0 43960 400
rect 44912 0 44968 400
rect 45920 0 45976 400
rect 46928 0 46984 400
rect 47936 0 47992 400
rect 48944 0 49000 400
rect 49952 0 50008 400
rect 50960 0 51016 400
rect 51968 0 52024 400
rect 52976 0 53032 400
rect 53984 0 54040 400
rect 54992 0 55048 400
rect 56000 0 56056 400
rect 57008 0 57064 400
rect 58016 0 58072 400
rect 59024 0 59080 400
rect 60032 0 60088 400
rect 61040 0 61096 400
rect 62048 0 62104 400
rect 63056 0 63112 400
rect 64064 0 64120 400
rect 65072 0 65128 400
rect 66080 0 66136 400
rect 67088 0 67144 400
rect 68096 0 68152 400
rect 69104 0 69160 400
rect 70112 0 70168 400
rect 71120 0 71176 400
rect 72128 0 72184 400
rect 73136 0 73192 400
rect 74144 0 74200 400
rect 75152 0 75208 400
rect 76160 0 76216 400
rect 77168 0 77224 400
rect 78176 0 78232 400
rect 79184 0 79240 400
rect 80192 0 80248 400
rect 81200 0 81256 400
rect 82208 0 82264 400
rect 83216 0 83272 400
rect 84224 0 84280 400
rect 85232 0 85288 400
rect 86240 0 86296 400
rect 87248 0 87304 400
rect 88256 0 88312 400
rect 89264 0 89320 400
rect 90272 0 90328 400
rect 91280 0 91336 400
rect 92288 0 92344 400
rect 93296 0 93352 400
rect 94304 0 94360 400
rect 95312 0 95368 400
rect 96320 0 96376 400
rect 97328 0 97384 400
rect 98336 0 98392 400
rect 99344 0 99400 400
rect 100352 0 100408 400
rect 101360 0 101416 400
rect 102368 0 102424 400
rect 103376 0 103432 400
<< obsm2 >>
rect 758 69570 1986 69650
rect 2102 69570 3330 69650
rect 3446 69570 4674 69650
rect 4790 69570 6018 69650
rect 6134 69570 7362 69650
rect 7478 69570 8706 69650
rect 8822 69570 10050 69650
rect 10166 69570 11394 69650
rect 11510 69570 12738 69650
rect 12854 69570 14082 69650
rect 14198 69570 15426 69650
rect 15542 69570 16770 69650
rect 16886 69570 18114 69650
rect 18230 69570 19458 69650
rect 19574 69570 20802 69650
rect 20918 69570 22146 69650
rect 22262 69570 23490 69650
rect 23606 69570 24834 69650
rect 24950 69570 26178 69650
rect 26294 69570 27522 69650
rect 27638 69570 28866 69650
rect 28982 69570 30210 69650
rect 30326 69570 31554 69650
rect 31670 69570 32898 69650
rect 33014 69570 34242 69650
rect 34358 69570 35586 69650
rect 35702 69570 36930 69650
rect 37046 69570 38274 69650
rect 38390 69570 39618 69650
rect 39734 69570 40962 69650
rect 41078 69570 42306 69650
rect 42422 69570 43650 69650
rect 43766 69570 44994 69650
rect 45110 69570 46338 69650
rect 46454 69570 47682 69650
rect 47798 69570 49026 69650
rect 49142 69570 50370 69650
rect 50486 69570 51714 69650
rect 51830 69570 53058 69650
rect 53174 69570 54402 69650
rect 54518 69570 55746 69650
rect 55862 69570 57090 69650
rect 57206 69570 58434 69650
rect 58550 69570 59778 69650
rect 59894 69570 61122 69650
rect 61238 69570 62466 69650
rect 62582 69570 63810 69650
rect 63926 69570 65154 69650
rect 65270 69570 66498 69650
rect 66614 69570 67842 69650
rect 67958 69570 69186 69650
rect 69302 69570 70530 69650
rect 70646 69570 71874 69650
rect 71990 69570 73218 69650
rect 73334 69570 74562 69650
rect 74678 69570 75906 69650
rect 76022 69570 77250 69650
rect 77366 69570 78594 69650
rect 78710 69570 79938 69650
rect 80054 69570 81282 69650
rect 81398 69570 82626 69650
rect 82742 69570 83970 69650
rect 84086 69570 85314 69650
rect 85430 69570 86658 69650
rect 86774 69570 88002 69650
rect 88118 69570 89346 69650
rect 89462 69570 90690 69650
rect 90806 69570 92034 69650
rect 92150 69570 93378 69650
rect 93494 69570 94722 69650
rect 94838 69570 96066 69650
rect 96182 69570 97410 69650
rect 97526 69570 98754 69650
rect 98870 69570 100098 69650
rect 100214 69570 101442 69650
rect 101558 69570 102786 69650
rect 102902 69570 104130 69650
rect 104246 69570 104370 69650
rect 686 430 104370 69570
rect 686 350 1538 430
rect 1654 350 2546 430
rect 2662 350 3554 430
rect 3670 350 4562 430
rect 4678 350 5570 430
rect 5686 350 6578 430
rect 6694 350 7586 430
rect 7702 350 8594 430
rect 8710 350 9602 430
rect 9718 350 10610 430
rect 10726 350 11618 430
rect 11734 350 12626 430
rect 12742 350 13634 430
rect 13750 350 14642 430
rect 14758 350 15650 430
rect 15766 350 16658 430
rect 16774 350 17666 430
rect 17782 350 18674 430
rect 18790 350 19682 430
rect 19798 350 20690 430
rect 20806 350 21698 430
rect 21814 350 22706 430
rect 22822 350 23714 430
rect 23830 350 24722 430
rect 24838 350 25730 430
rect 25846 350 26738 430
rect 26854 350 27746 430
rect 27862 350 28754 430
rect 28870 350 29762 430
rect 29878 350 30770 430
rect 30886 350 31778 430
rect 31894 350 32786 430
rect 32902 350 33794 430
rect 33910 350 34802 430
rect 34918 350 35810 430
rect 35926 350 36818 430
rect 36934 350 37826 430
rect 37942 350 38834 430
rect 38950 350 39842 430
rect 39958 350 40850 430
rect 40966 350 41858 430
rect 41974 350 42866 430
rect 42982 350 43874 430
rect 43990 350 44882 430
rect 44998 350 45890 430
rect 46006 350 46898 430
rect 47014 350 47906 430
rect 48022 350 48914 430
rect 49030 350 49922 430
rect 50038 350 50930 430
rect 51046 350 51938 430
rect 52054 350 52946 430
rect 53062 350 53954 430
rect 54070 350 54962 430
rect 55078 350 55970 430
rect 56086 350 56978 430
rect 57094 350 57986 430
rect 58102 350 58994 430
rect 59110 350 60002 430
rect 60118 350 61010 430
rect 61126 350 62018 430
rect 62134 350 63026 430
rect 63142 350 64034 430
rect 64150 350 65042 430
rect 65158 350 66050 430
rect 66166 350 67058 430
rect 67174 350 68066 430
rect 68182 350 69074 430
rect 69190 350 70082 430
rect 70198 350 71090 430
rect 71206 350 72098 430
rect 72214 350 73106 430
rect 73222 350 74114 430
rect 74230 350 75122 430
rect 75238 350 76130 430
rect 76246 350 77138 430
rect 77254 350 78146 430
rect 78262 350 79154 430
rect 79270 350 80162 430
rect 80278 350 81170 430
rect 81286 350 82178 430
rect 82294 350 83186 430
rect 83302 350 84194 430
rect 84310 350 85202 430
rect 85318 350 86210 430
rect 86326 350 87218 430
rect 87334 350 88226 430
rect 88342 350 89234 430
rect 89350 350 90242 430
rect 90358 350 91250 430
rect 91366 350 92258 430
rect 92374 350 93266 430
rect 93382 350 94274 430
rect 94390 350 95282 430
rect 95398 350 96290 430
rect 96406 350 97298 430
rect 97414 350 98306 430
rect 98422 350 99314 430
rect 99430 350 100322 430
rect 100438 350 101330 430
rect 101446 350 102338 430
rect 102454 350 103346 430
rect 103462 350 104370 430
<< metal3 >>
rect 0 67872 400 67928
rect 0 67200 400 67256
rect 0 66528 400 66584
rect 104600 66192 105000 66248
rect 0 65856 400 65912
rect 104600 65520 105000 65576
rect 0 65184 400 65240
rect 104600 64848 105000 64904
rect 0 64512 400 64568
rect 104600 64176 105000 64232
rect 0 63840 400 63896
rect 104600 63504 105000 63560
rect 0 63168 400 63224
rect 104600 62832 105000 62888
rect 0 62496 400 62552
rect 104600 62160 105000 62216
rect 0 61824 400 61880
rect 104600 61488 105000 61544
rect 0 61152 400 61208
rect 104600 60816 105000 60872
rect 0 60480 400 60536
rect 104600 60144 105000 60200
rect 0 59808 400 59864
rect 104600 59472 105000 59528
rect 0 59136 400 59192
rect 104600 58800 105000 58856
rect 0 58464 400 58520
rect 104600 58128 105000 58184
rect 0 57792 400 57848
rect 104600 57456 105000 57512
rect 0 57120 400 57176
rect 104600 56784 105000 56840
rect 0 56448 400 56504
rect 104600 56112 105000 56168
rect 0 55776 400 55832
rect 104600 55440 105000 55496
rect 0 55104 400 55160
rect 104600 54768 105000 54824
rect 0 54432 400 54488
rect 104600 54096 105000 54152
rect 0 53760 400 53816
rect 104600 53424 105000 53480
rect 0 53088 400 53144
rect 104600 52752 105000 52808
rect 0 52416 400 52472
rect 104600 52080 105000 52136
rect 0 51744 400 51800
rect 104600 51408 105000 51464
rect 0 51072 400 51128
rect 104600 50736 105000 50792
rect 0 50400 400 50456
rect 104600 50064 105000 50120
rect 0 49728 400 49784
rect 104600 49392 105000 49448
rect 0 49056 400 49112
rect 104600 48720 105000 48776
rect 0 48384 400 48440
rect 104600 48048 105000 48104
rect 0 47712 400 47768
rect 104600 47376 105000 47432
rect 0 47040 400 47096
rect 104600 46704 105000 46760
rect 0 46368 400 46424
rect 104600 46032 105000 46088
rect 0 45696 400 45752
rect 104600 45360 105000 45416
rect 0 45024 400 45080
rect 104600 44688 105000 44744
rect 0 44352 400 44408
rect 104600 44016 105000 44072
rect 0 43680 400 43736
rect 104600 43344 105000 43400
rect 0 43008 400 43064
rect 104600 42672 105000 42728
rect 0 42336 400 42392
rect 104600 42000 105000 42056
rect 0 41664 400 41720
rect 104600 41328 105000 41384
rect 0 40992 400 41048
rect 104600 40656 105000 40712
rect 0 40320 400 40376
rect 104600 39984 105000 40040
rect 0 39648 400 39704
rect 104600 39312 105000 39368
rect 0 38976 400 39032
rect 104600 38640 105000 38696
rect 0 38304 400 38360
rect 104600 37968 105000 38024
rect 0 37632 400 37688
rect 104600 37296 105000 37352
rect 0 36960 400 37016
rect 104600 36624 105000 36680
rect 0 36288 400 36344
rect 104600 35952 105000 36008
rect 0 35616 400 35672
rect 104600 35280 105000 35336
rect 0 34944 400 35000
rect 104600 34608 105000 34664
rect 0 34272 400 34328
rect 104600 33936 105000 33992
rect 0 33600 400 33656
rect 104600 33264 105000 33320
rect 0 32928 400 32984
rect 104600 32592 105000 32648
rect 0 32256 400 32312
rect 104600 31920 105000 31976
rect 0 31584 400 31640
rect 104600 31248 105000 31304
rect 0 30912 400 30968
rect 104600 30576 105000 30632
rect 0 30240 400 30296
rect 104600 29904 105000 29960
rect 0 29568 400 29624
rect 104600 29232 105000 29288
rect 0 28896 400 28952
rect 104600 28560 105000 28616
rect 0 28224 400 28280
rect 104600 27888 105000 27944
rect 0 27552 400 27608
rect 104600 27216 105000 27272
rect 0 26880 400 26936
rect 104600 26544 105000 26600
rect 0 26208 400 26264
rect 104600 25872 105000 25928
rect 0 25536 400 25592
rect 104600 25200 105000 25256
rect 0 24864 400 24920
rect 104600 24528 105000 24584
rect 0 24192 400 24248
rect 104600 23856 105000 23912
rect 0 23520 400 23576
rect 104600 23184 105000 23240
rect 0 22848 400 22904
rect 104600 22512 105000 22568
rect 0 22176 400 22232
rect 104600 21840 105000 21896
rect 0 21504 400 21560
rect 104600 21168 105000 21224
rect 0 20832 400 20888
rect 104600 20496 105000 20552
rect 0 20160 400 20216
rect 104600 19824 105000 19880
rect 0 19488 400 19544
rect 104600 19152 105000 19208
rect 0 18816 400 18872
rect 104600 18480 105000 18536
rect 0 18144 400 18200
rect 104600 17808 105000 17864
rect 0 17472 400 17528
rect 104600 17136 105000 17192
rect 0 16800 400 16856
rect 104600 16464 105000 16520
rect 0 16128 400 16184
rect 104600 15792 105000 15848
rect 0 15456 400 15512
rect 104600 15120 105000 15176
rect 0 14784 400 14840
rect 104600 14448 105000 14504
rect 0 14112 400 14168
rect 104600 13776 105000 13832
rect 0 13440 400 13496
rect 104600 13104 105000 13160
rect 0 12768 400 12824
rect 104600 12432 105000 12488
rect 0 12096 400 12152
rect 104600 11760 105000 11816
rect 0 11424 400 11480
rect 104600 11088 105000 11144
rect 0 10752 400 10808
rect 104600 10416 105000 10472
rect 0 10080 400 10136
rect 104600 9744 105000 9800
rect 0 9408 400 9464
rect 104600 9072 105000 9128
rect 0 8736 400 8792
rect 104600 8400 105000 8456
rect 0 8064 400 8120
rect 104600 7728 105000 7784
rect 0 7392 400 7448
rect 104600 7056 105000 7112
rect 0 6720 400 6776
rect 104600 6384 105000 6440
rect 0 6048 400 6104
rect 104600 5712 105000 5768
rect 0 5376 400 5432
rect 104600 5040 105000 5096
rect 0 4704 400 4760
rect 104600 4368 105000 4424
rect 0 4032 400 4088
rect 104600 3696 105000 3752
rect 0 3360 400 3416
rect 0 2688 400 2744
rect 0 2016 400 2072
<< obsm3 >>
rect 400 67958 104650 68474
rect 430 67842 104650 67958
rect 400 67286 104650 67842
rect 430 67170 104650 67286
rect 400 66614 104650 67170
rect 430 66498 104650 66614
rect 400 66278 104650 66498
rect 400 66162 104570 66278
rect 400 65942 104650 66162
rect 430 65826 104650 65942
rect 400 65606 104650 65826
rect 400 65490 104570 65606
rect 400 65270 104650 65490
rect 430 65154 104650 65270
rect 400 64934 104650 65154
rect 400 64818 104570 64934
rect 400 64598 104650 64818
rect 430 64482 104650 64598
rect 400 64262 104650 64482
rect 400 64146 104570 64262
rect 400 63926 104650 64146
rect 430 63810 104650 63926
rect 400 63590 104650 63810
rect 400 63474 104570 63590
rect 400 63254 104650 63474
rect 430 63138 104650 63254
rect 400 62918 104650 63138
rect 400 62802 104570 62918
rect 400 62582 104650 62802
rect 430 62466 104650 62582
rect 400 62246 104650 62466
rect 400 62130 104570 62246
rect 400 61910 104650 62130
rect 430 61794 104650 61910
rect 400 61574 104650 61794
rect 400 61458 104570 61574
rect 400 61238 104650 61458
rect 430 61122 104650 61238
rect 400 60902 104650 61122
rect 400 60786 104570 60902
rect 400 60566 104650 60786
rect 430 60450 104650 60566
rect 400 60230 104650 60450
rect 400 60114 104570 60230
rect 400 59894 104650 60114
rect 430 59778 104650 59894
rect 400 59558 104650 59778
rect 400 59442 104570 59558
rect 400 59222 104650 59442
rect 430 59106 104650 59222
rect 400 58886 104650 59106
rect 400 58770 104570 58886
rect 400 58550 104650 58770
rect 430 58434 104650 58550
rect 400 58214 104650 58434
rect 400 58098 104570 58214
rect 400 57878 104650 58098
rect 430 57762 104650 57878
rect 400 57542 104650 57762
rect 400 57426 104570 57542
rect 400 57206 104650 57426
rect 430 57090 104650 57206
rect 400 56870 104650 57090
rect 400 56754 104570 56870
rect 400 56534 104650 56754
rect 430 56418 104650 56534
rect 400 56198 104650 56418
rect 400 56082 104570 56198
rect 400 55862 104650 56082
rect 430 55746 104650 55862
rect 400 55526 104650 55746
rect 400 55410 104570 55526
rect 400 55190 104650 55410
rect 430 55074 104650 55190
rect 400 54854 104650 55074
rect 400 54738 104570 54854
rect 400 54518 104650 54738
rect 430 54402 104650 54518
rect 400 54182 104650 54402
rect 400 54066 104570 54182
rect 400 53846 104650 54066
rect 430 53730 104650 53846
rect 400 53510 104650 53730
rect 400 53394 104570 53510
rect 400 53174 104650 53394
rect 430 53058 104650 53174
rect 400 52838 104650 53058
rect 400 52722 104570 52838
rect 400 52502 104650 52722
rect 430 52386 104650 52502
rect 400 52166 104650 52386
rect 400 52050 104570 52166
rect 400 51830 104650 52050
rect 430 51714 104650 51830
rect 400 51494 104650 51714
rect 400 51378 104570 51494
rect 400 51158 104650 51378
rect 430 51042 104650 51158
rect 400 50822 104650 51042
rect 400 50706 104570 50822
rect 400 50486 104650 50706
rect 430 50370 104650 50486
rect 400 50150 104650 50370
rect 400 50034 104570 50150
rect 400 49814 104650 50034
rect 430 49698 104650 49814
rect 400 49478 104650 49698
rect 400 49362 104570 49478
rect 400 49142 104650 49362
rect 430 49026 104650 49142
rect 400 48806 104650 49026
rect 400 48690 104570 48806
rect 400 48470 104650 48690
rect 430 48354 104650 48470
rect 400 48134 104650 48354
rect 400 48018 104570 48134
rect 400 47798 104650 48018
rect 430 47682 104650 47798
rect 400 47462 104650 47682
rect 400 47346 104570 47462
rect 400 47126 104650 47346
rect 430 47010 104650 47126
rect 400 46790 104650 47010
rect 400 46674 104570 46790
rect 400 46454 104650 46674
rect 430 46338 104650 46454
rect 400 46118 104650 46338
rect 400 46002 104570 46118
rect 400 45782 104650 46002
rect 430 45666 104650 45782
rect 400 45446 104650 45666
rect 400 45330 104570 45446
rect 400 45110 104650 45330
rect 430 44994 104650 45110
rect 400 44774 104650 44994
rect 400 44658 104570 44774
rect 400 44438 104650 44658
rect 430 44322 104650 44438
rect 400 44102 104650 44322
rect 400 43986 104570 44102
rect 400 43766 104650 43986
rect 430 43650 104650 43766
rect 400 43430 104650 43650
rect 400 43314 104570 43430
rect 400 43094 104650 43314
rect 430 42978 104650 43094
rect 400 42758 104650 42978
rect 400 42642 104570 42758
rect 400 42422 104650 42642
rect 430 42306 104650 42422
rect 400 42086 104650 42306
rect 400 41970 104570 42086
rect 400 41750 104650 41970
rect 430 41634 104650 41750
rect 400 41414 104650 41634
rect 400 41298 104570 41414
rect 400 41078 104650 41298
rect 430 40962 104650 41078
rect 400 40742 104650 40962
rect 400 40626 104570 40742
rect 400 40406 104650 40626
rect 430 40290 104650 40406
rect 400 40070 104650 40290
rect 400 39954 104570 40070
rect 400 39734 104650 39954
rect 430 39618 104650 39734
rect 400 39398 104650 39618
rect 400 39282 104570 39398
rect 400 39062 104650 39282
rect 430 38946 104650 39062
rect 400 38726 104650 38946
rect 400 38610 104570 38726
rect 400 38390 104650 38610
rect 430 38274 104650 38390
rect 400 38054 104650 38274
rect 400 37938 104570 38054
rect 400 37718 104650 37938
rect 430 37602 104650 37718
rect 400 37382 104650 37602
rect 400 37266 104570 37382
rect 400 37046 104650 37266
rect 430 36930 104650 37046
rect 400 36710 104650 36930
rect 400 36594 104570 36710
rect 400 36374 104650 36594
rect 430 36258 104650 36374
rect 400 36038 104650 36258
rect 400 35922 104570 36038
rect 400 35702 104650 35922
rect 430 35586 104650 35702
rect 400 35366 104650 35586
rect 400 35250 104570 35366
rect 400 35030 104650 35250
rect 430 34914 104650 35030
rect 400 34694 104650 34914
rect 400 34578 104570 34694
rect 400 34358 104650 34578
rect 430 34242 104650 34358
rect 400 34022 104650 34242
rect 400 33906 104570 34022
rect 400 33686 104650 33906
rect 430 33570 104650 33686
rect 400 33350 104650 33570
rect 400 33234 104570 33350
rect 400 33014 104650 33234
rect 430 32898 104650 33014
rect 400 32678 104650 32898
rect 400 32562 104570 32678
rect 400 32342 104650 32562
rect 430 32226 104650 32342
rect 400 32006 104650 32226
rect 400 31890 104570 32006
rect 400 31670 104650 31890
rect 430 31554 104650 31670
rect 400 31334 104650 31554
rect 400 31218 104570 31334
rect 400 30998 104650 31218
rect 430 30882 104650 30998
rect 400 30662 104650 30882
rect 400 30546 104570 30662
rect 400 30326 104650 30546
rect 430 30210 104650 30326
rect 400 29990 104650 30210
rect 400 29874 104570 29990
rect 400 29654 104650 29874
rect 430 29538 104650 29654
rect 400 29318 104650 29538
rect 400 29202 104570 29318
rect 400 28982 104650 29202
rect 430 28866 104650 28982
rect 400 28646 104650 28866
rect 400 28530 104570 28646
rect 400 28310 104650 28530
rect 430 28194 104650 28310
rect 400 27974 104650 28194
rect 400 27858 104570 27974
rect 400 27638 104650 27858
rect 430 27522 104650 27638
rect 400 27302 104650 27522
rect 400 27186 104570 27302
rect 400 26966 104650 27186
rect 430 26850 104650 26966
rect 400 26630 104650 26850
rect 400 26514 104570 26630
rect 400 26294 104650 26514
rect 430 26178 104650 26294
rect 400 25958 104650 26178
rect 400 25842 104570 25958
rect 400 25622 104650 25842
rect 430 25506 104650 25622
rect 400 25286 104650 25506
rect 400 25170 104570 25286
rect 400 24950 104650 25170
rect 430 24834 104650 24950
rect 400 24614 104650 24834
rect 400 24498 104570 24614
rect 400 24278 104650 24498
rect 430 24162 104650 24278
rect 400 23942 104650 24162
rect 400 23826 104570 23942
rect 400 23606 104650 23826
rect 430 23490 104650 23606
rect 400 23270 104650 23490
rect 400 23154 104570 23270
rect 400 22934 104650 23154
rect 430 22818 104650 22934
rect 400 22598 104650 22818
rect 400 22482 104570 22598
rect 400 22262 104650 22482
rect 430 22146 104650 22262
rect 400 21926 104650 22146
rect 400 21810 104570 21926
rect 400 21590 104650 21810
rect 430 21474 104650 21590
rect 400 21254 104650 21474
rect 400 21138 104570 21254
rect 400 20918 104650 21138
rect 430 20802 104650 20918
rect 400 20582 104650 20802
rect 400 20466 104570 20582
rect 400 20246 104650 20466
rect 430 20130 104650 20246
rect 400 19910 104650 20130
rect 400 19794 104570 19910
rect 400 19574 104650 19794
rect 430 19458 104650 19574
rect 400 19238 104650 19458
rect 400 19122 104570 19238
rect 400 18902 104650 19122
rect 430 18786 104650 18902
rect 400 18566 104650 18786
rect 400 18450 104570 18566
rect 400 18230 104650 18450
rect 430 18114 104650 18230
rect 400 17894 104650 18114
rect 400 17778 104570 17894
rect 400 17558 104650 17778
rect 430 17442 104650 17558
rect 400 17222 104650 17442
rect 400 17106 104570 17222
rect 400 16886 104650 17106
rect 430 16770 104650 16886
rect 400 16550 104650 16770
rect 400 16434 104570 16550
rect 400 16214 104650 16434
rect 430 16098 104650 16214
rect 400 15878 104650 16098
rect 400 15762 104570 15878
rect 400 15542 104650 15762
rect 430 15426 104650 15542
rect 400 15206 104650 15426
rect 400 15090 104570 15206
rect 400 14870 104650 15090
rect 430 14754 104650 14870
rect 400 14534 104650 14754
rect 400 14418 104570 14534
rect 400 14198 104650 14418
rect 430 14082 104650 14198
rect 400 13862 104650 14082
rect 400 13746 104570 13862
rect 400 13526 104650 13746
rect 430 13410 104650 13526
rect 400 13190 104650 13410
rect 400 13074 104570 13190
rect 400 12854 104650 13074
rect 430 12738 104650 12854
rect 400 12518 104650 12738
rect 400 12402 104570 12518
rect 400 12182 104650 12402
rect 430 12066 104650 12182
rect 400 11846 104650 12066
rect 400 11730 104570 11846
rect 400 11510 104650 11730
rect 430 11394 104650 11510
rect 400 11174 104650 11394
rect 400 11058 104570 11174
rect 400 10838 104650 11058
rect 430 10722 104650 10838
rect 400 10502 104650 10722
rect 400 10386 104570 10502
rect 400 10166 104650 10386
rect 430 10050 104650 10166
rect 400 9830 104650 10050
rect 400 9714 104570 9830
rect 400 9494 104650 9714
rect 430 9378 104650 9494
rect 400 9158 104650 9378
rect 400 9042 104570 9158
rect 400 8822 104650 9042
rect 430 8706 104650 8822
rect 400 8486 104650 8706
rect 400 8370 104570 8486
rect 400 8150 104650 8370
rect 430 8034 104650 8150
rect 400 7814 104650 8034
rect 400 7698 104570 7814
rect 400 7478 104650 7698
rect 430 7362 104650 7478
rect 400 7142 104650 7362
rect 400 7026 104570 7142
rect 400 6806 104650 7026
rect 430 6690 104650 6806
rect 400 6470 104650 6690
rect 400 6354 104570 6470
rect 400 6134 104650 6354
rect 430 6018 104650 6134
rect 400 5798 104650 6018
rect 400 5682 104570 5798
rect 400 5462 104650 5682
rect 430 5346 104650 5462
rect 400 5126 104650 5346
rect 400 5010 104570 5126
rect 400 4790 104650 5010
rect 430 4674 104650 4790
rect 400 4454 104650 4674
rect 400 4338 104570 4454
rect 400 4118 104650 4338
rect 430 4002 104650 4118
rect 400 3782 104650 4002
rect 400 3666 104570 3782
rect 400 3446 104650 3666
rect 430 3330 104650 3446
rect 400 2774 104650 3330
rect 430 2658 104650 2774
rect 400 2102 104650 2658
rect 430 1986 104650 2102
rect 400 1414 104650 1986
<< metal4 >>
rect 2224 1538 2384 68238
rect 9904 1538 10064 68238
rect 17584 1538 17744 68238
rect 25264 1538 25424 68238
rect 32944 1538 33104 68238
rect 40624 1538 40784 68238
rect 48304 1538 48464 68238
rect 55984 1538 56144 68238
rect 63664 1538 63824 68238
rect 71344 1538 71504 68238
rect 79024 1538 79184 68238
rect 86704 1538 86864 68238
rect 94384 1538 94544 68238
rect 102064 1538 102224 68238
<< obsm4 >>
rect 13062 6001 17554 66575
rect 17774 6001 25234 66575
rect 25454 6001 32914 66575
rect 33134 6001 40594 66575
rect 40814 6001 48274 66575
rect 48494 6001 55954 66575
rect 56174 6001 63634 66575
rect 63854 6001 71314 66575
rect 71534 6001 78994 66575
rect 79214 6001 86674 66575
rect 86894 6001 94354 66575
rect 94574 6001 99890 66575
<< labels >>
rlabel metal3 s 0 40992 400 41048 6 RAM_end_addr[0]
port 1 nsew signal output
rlabel metal3 s 0 47712 400 47768 6 RAM_end_addr[10]
port 2 nsew signal output
rlabel metal3 s 0 48384 400 48440 6 RAM_end_addr[11]
port 3 nsew signal output
rlabel metal3 s 0 49056 400 49112 6 RAM_end_addr[12]
port 4 nsew signal output
rlabel metal3 s 0 49728 400 49784 6 RAM_end_addr[13]
port 5 nsew signal output
rlabel metal3 s 0 50400 400 50456 6 RAM_end_addr[14]
port 6 nsew signal output
rlabel metal3 s 0 51072 400 51128 6 RAM_end_addr[15]
port 7 nsew signal output
rlabel metal3 s 0 41664 400 41720 6 RAM_end_addr[1]
port 8 nsew signal output
rlabel metal3 s 0 42336 400 42392 6 RAM_end_addr[2]
port 9 nsew signal output
rlabel metal3 s 0 43008 400 43064 6 RAM_end_addr[3]
port 10 nsew signal output
rlabel metal3 s 0 43680 400 43736 6 RAM_end_addr[4]
port 11 nsew signal output
rlabel metal3 s 0 44352 400 44408 6 RAM_end_addr[5]
port 12 nsew signal output
rlabel metal3 s 0 45024 400 45080 6 RAM_end_addr[6]
port 13 nsew signal output
rlabel metal3 s 0 45696 400 45752 6 RAM_end_addr[7]
port 14 nsew signal output
rlabel metal3 s 0 46368 400 46424 6 RAM_end_addr[8]
port 15 nsew signal output
rlabel metal3 s 0 47040 400 47096 6 RAM_end_addr[9]
port 16 nsew signal output
rlabel metal3 s 0 27552 400 27608 6 RAM_start_addr[0]
port 17 nsew signal output
rlabel metal3 s 0 34272 400 34328 6 RAM_start_addr[10]
port 18 nsew signal output
rlabel metal3 s 0 34944 400 35000 6 RAM_start_addr[11]
port 19 nsew signal output
rlabel metal3 s 0 35616 400 35672 6 RAM_start_addr[12]
port 20 nsew signal output
rlabel metal3 s 0 36288 400 36344 6 RAM_start_addr[13]
port 21 nsew signal output
rlabel metal3 s 0 36960 400 37016 6 RAM_start_addr[14]
port 22 nsew signal output
rlabel metal3 s 0 37632 400 37688 6 RAM_start_addr[15]
port 23 nsew signal output
rlabel metal3 s 0 28224 400 28280 6 RAM_start_addr[1]
port 24 nsew signal output
rlabel metal3 s 0 28896 400 28952 6 RAM_start_addr[2]
port 25 nsew signal output
rlabel metal3 s 0 29568 400 29624 6 RAM_start_addr[3]
port 26 nsew signal output
rlabel metal3 s 0 30240 400 30296 6 RAM_start_addr[4]
port 27 nsew signal output
rlabel metal3 s 0 30912 400 30968 6 RAM_start_addr[5]
port 28 nsew signal output
rlabel metal3 s 0 31584 400 31640 6 RAM_start_addr[6]
port 29 nsew signal output
rlabel metal3 s 0 32256 400 32312 6 RAM_start_addr[7]
port 30 nsew signal output
rlabel metal3 s 0 32928 400 32984 6 RAM_start_addr[8]
port 31 nsew signal output
rlabel metal3 s 0 33600 400 33656 6 RAM_start_addr[9]
port 32 nsew signal output
rlabel metal2 s 66528 69600 66584 70000 6 WEb_ram
port 33 nsew signal output
rlabel metal3 s 0 40320 400 40376 6 boot_rom_en
port 34 nsew signal output
rlabel metal2 s 47712 69600 47768 70000 6 bus_addr[0]
port 35 nsew signal output
rlabel metal2 s 49056 69600 49112 70000 6 bus_addr[1]
port 36 nsew signal output
rlabel metal2 s 50400 69600 50456 70000 6 bus_addr[2]
port 37 nsew signal output
rlabel metal2 s 51744 69600 51800 70000 6 bus_addr[3]
port 38 nsew signal output
rlabel metal2 s 53088 69600 53144 70000 6 bus_addr[4]
port 39 nsew signal output
rlabel metal2 s 54432 69600 54488 70000 6 bus_addr[5]
port 40 nsew signal output
rlabel metal2 s 46368 69600 46424 70000 6 bus_cyc
port 41 nsew signal output
rlabel metal2 s 35616 69600 35672 70000 6 bus_data_out[0]
port 42 nsew signal output
rlabel metal2 s 36960 69600 37016 70000 6 bus_data_out[1]
port 43 nsew signal output
rlabel metal2 s 38304 69600 38360 70000 6 bus_data_out[2]
port 44 nsew signal output
rlabel metal2 s 39648 69600 39704 70000 6 bus_data_out[3]
port 45 nsew signal output
rlabel metal2 s 40992 69600 41048 70000 6 bus_data_out[4]
port 46 nsew signal output
rlabel metal2 s 42336 69600 42392 70000 6 bus_data_out[5]
port 47 nsew signal output
rlabel metal2 s 43680 69600 43736 70000 6 bus_data_out[6]
port 48 nsew signal output
rlabel metal2 s 45024 69600 45080 70000 6 bus_data_out[7]
port 49 nsew signal output
rlabel metal3 s 104600 44016 105000 44072 6 bus_in_gpios[0]
port 50 nsew signal input
rlabel metal3 s 104600 44688 105000 44744 6 bus_in_gpios[1]
port 51 nsew signal input
rlabel metal3 s 104600 45360 105000 45416 6 bus_in_gpios[2]
port 52 nsew signal input
rlabel metal3 s 104600 46032 105000 46088 6 bus_in_gpios[3]
port 53 nsew signal input
rlabel metal3 s 104600 46704 105000 46760 6 bus_in_gpios[4]
port 54 nsew signal input
rlabel metal3 s 104600 47376 105000 47432 6 bus_in_gpios[5]
port 55 nsew signal input
rlabel metal3 s 104600 48048 105000 48104 6 bus_in_gpios[6]
port 56 nsew signal input
rlabel metal3 s 104600 48720 105000 48776 6 bus_in_gpios[7]
port 57 nsew signal input
rlabel metal2 s 55776 69600 55832 70000 6 bus_in_serial_ports[0]
port 58 nsew signal input
rlabel metal2 s 57120 69600 57176 70000 6 bus_in_serial_ports[1]
port 59 nsew signal input
rlabel metal2 s 58464 69600 58520 70000 6 bus_in_serial_ports[2]
port 60 nsew signal input
rlabel metal2 s 59808 69600 59864 70000 6 bus_in_serial_ports[3]
port 61 nsew signal input
rlabel metal2 s 61152 69600 61208 70000 6 bus_in_serial_ports[4]
port 62 nsew signal input
rlabel metal2 s 62496 69600 62552 70000 6 bus_in_serial_ports[5]
port 63 nsew signal input
rlabel metal2 s 63840 69600 63896 70000 6 bus_in_serial_ports[6]
port 64 nsew signal input
rlabel metal2 s 65184 69600 65240 70000 6 bus_in_serial_ports[7]
port 65 nsew signal input
rlabel metal3 s 104600 50736 105000 50792 6 bus_in_sid[0]
port 66 nsew signal input
rlabel metal3 s 104600 51408 105000 51464 6 bus_in_sid[1]
port 67 nsew signal input
rlabel metal3 s 104600 52080 105000 52136 6 bus_in_sid[2]
port 68 nsew signal input
rlabel metal3 s 104600 52752 105000 52808 6 bus_in_sid[3]
port 69 nsew signal input
rlabel metal3 s 104600 53424 105000 53480 6 bus_in_sid[4]
port 70 nsew signal input
rlabel metal3 s 104600 54096 105000 54152 6 bus_in_sid[5]
port 71 nsew signal input
rlabel metal3 s 104600 54768 105000 54824 6 bus_in_sid[6]
port 72 nsew signal input
rlabel metal3 s 104600 55440 105000 55496 6 bus_in_sid[7]
port 73 nsew signal input
rlabel metal2 s 94752 69600 94808 70000 6 bus_in_timers[0]
port 74 nsew signal input
rlabel metal2 s 96096 69600 96152 70000 6 bus_in_timers[1]
port 75 nsew signal input
rlabel metal2 s 97440 69600 97496 70000 6 bus_in_timers[2]
port 76 nsew signal input
rlabel metal2 s 98784 69600 98840 70000 6 bus_in_timers[3]
port 77 nsew signal input
rlabel metal2 s 100128 69600 100184 70000 6 bus_in_timers[4]
port 78 nsew signal input
rlabel metal2 s 101472 69600 101528 70000 6 bus_in_timers[5]
port 79 nsew signal input
rlabel metal2 s 102816 69600 102872 70000 6 bus_in_timers[6]
port 80 nsew signal input
rlabel metal2 s 104160 69600 104216 70000 6 bus_in_timers[7]
port 81 nsew signal input
rlabel metal3 s 104600 43344 105000 43400 6 bus_we_gpios
port 82 nsew signal output
rlabel metal2 s 93408 69600 93464 70000 6 bus_we_serial_ports
port 83 nsew signal output
rlabel metal3 s 104600 50064 105000 50120 6 bus_we_sid
port 84 nsew signal output
rlabel metal2 s 92064 69600 92120 70000 6 bus_we_timers
port 85 nsew signal output
rlabel metal3 s 0 38304 400 38360 6 cs_port[0]
port 86 nsew signal output
rlabel metal3 s 0 38976 400 39032 6 cs_port[1]
port 87 nsew signal output
rlabel metal3 s 0 39648 400 39704 6 cs_port[2]
port 88 nsew signal output
rlabel metal2 s 672 69600 728 70000 6 io_in[0]
port 89 nsew signal input
rlabel metal2 s 14112 69600 14168 70000 6 io_in[10]
port 90 nsew signal input
rlabel metal2 s 15456 69600 15512 70000 6 io_in[11]
port 91 nsew signal input
rlabel metal2 s 16800 69600 16856 70000 6 io_in[12]
port 92 nsew signal input
rlabel metal2 s 18144 69600 18200 70000 6 io_in[13]
port 93 nsew signal input
rlabel metal2 s 19488 69600 19544 70000 6 io_in[14]
port 94 nsew signal input
rlabel metal2 s 20832 69600 20888 70000 6 io_in[15]
port 95 nsew signal input
rlabel metal2 s 22176 69600 22232 70000 6 io_in[16]
port 96 nsew signal input
rlabel metal2 s 23520 69600 23576 70000 6 io_in[17]
port 97 nsew signal input
rlabel metal2 s 24864 69600 24920 70000 6 io_in[18]
port 98 nsew signal input
rlabel metal2 s 2016 69600 2072 70000 6 io_in[1]
port 99 nsew signal input
rlabel metal2 s 3360 69600 3416 70000 6 io_in[2]
port 100 nsew signal input
rlabel metal2 s 4704 69600 4760 70000 6 io_in[3]
port 101 nsew signal input
rlabel metal2 s 6048 69600 6104 70000 6 io_in[4]
port 102 nsew signal input
rlabel metal2 s 7392 69600 7448 70000 6 io_in[5]
port 103 nsew signal input
rlabel metal2 s 8736 69600 8792 70000 6 io_in[6]
port 104 nsew signal input
rlabel metal2 s 10080 69600 10136 70000 6 io_in[7]
port 105 nsew signal input
rlabel metal2 s 11424 69600 11480 70000 6 io_in[8]
port 106 nsew signal input
rlabel metal2 s 12768 69600 12824 70000 6 io_in[9]
port 107 nsew signal input
rlabel metal3 s 0 14784 400 14840 6 io_oeb[0]
port 108 nsew signal output
rlabel metal3 s 0 21504 400 21560 6 io_oeb[10]
port 109 nsew signal output
rlabel metal3 s 0 22176 400 22232 6 io_oeb[11]
port 110 nsew signal output
rlabel metal3 s 0 22848 400 22904 6 io_oeb[12]
port 111 nsew signal output
rlabel metal3 s 0 23520 400 23576 6 io_oeb[13]
port 112 nsew signal output
rlabel metal3 s 0 24192 400 24248 6 io_oeb[14]
port 113 nsew signal output
rlabel metal3 s 0 24864 400 24920 6 io_oeb[15]
port 114 nsew signal output
rlabel metal3 s 0 25536 400 25592 6 io_oeb[16]
port 115 nsew signal output
rlabel metal3 s 0 26208 400 26264 6 io_oeb[17]
port 116 nsew signal output
rlabel metal3 s 0 26880 400 26936 6 io_oeb[18]
port 117 nsew signal output
rlabel metal3 s 0 15456 400 15512 6 io_oeb[1]
port 118 nsew signal output
rlabel metal3 s 0 16128 400 16184 6 io_oeb[2]
port 119 nsew signal output
rlabel metal3 s 0 16800 400 16856 6 io_oeb[3]
port 120 nsew signal output
rlabel metal3 s 0 17472 400 17528 6 io_oeb[4]
port 121 nsew signal output
rlabel metal3 s 0 18144 400 18200 6 io_oeb[5]
port 122 nsew signal output
rlabel metal3 s 0 18816 400 18872 6 io_oeb[6]
port 123 nsew signal output
rlabel metal3 s 0 19488 400 19544 6 io_oeb[7]
port 124 nsew signal output
rlabel metal3 s 0 20160 400 20216 6 io_oeb[8]
port 125 nsew signal output
rlabel metal3 s 0 20832 400 20888 6 io_oeb[9]
port 126 nsew signal output
rlabel metal3 s 0 2016 400 2072 6 io_out[0]
port 127 nsew signal output
rlabel metal3 s 0 8736 400 8792 6 io_out[10]
port 128 nsew signal output
rlabel metal3 s 0 9408 400 9464 6 io_out[11]
port 129 nsew signal output
rlabel metal3 s 0 10080 400 10136 6 io_out[12]
port 130 nsew signal output
rlabel metal3 s 0 10752 400 10808 6 io_out[13]
port 131 nsew signal output
rlabel metal3 s 0 11424 400 11480 6 io_out[14]
port 132 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 io_out[15]
port 133 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 io_out[16]
port 134 nsew signal output
rlabel metal3 s 0 13440 400 13496 6 io_out[17]
port 135 nsew signal output
rlabel metal3 s 0 14112 400 14168 6 io_out[18]
port 136 nsew signal output
rlabel metal3 s 0 2688 400 2744 6 io_out[1]
port 137 nsew signal output
rlabel metal3 s 0 3360 400 3416 6 io_out[2]
port 138 nsew signal output
rlabel metal3 s 0 4032 400 4088 6 io_out[3]
port 139 nsew signal output
rlabel metal3 s 0 4704 400 4760 6 io_out[4]
port 140 nsew signal output
rlabel metal3 s 0 5376 400 5432 6 io_out[5]
port 141 nsew signal output
rlabel metal3 s 0 6048 400 6104 6 io_out[6]
port 142 nsew signal output
rlabel metal3 s 0 6720 400 6776 6 io_out[7]
port 143 nsew signal output
rlabel metal3 s 0 7392 400 7448 6 io_out[8]
port 144 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 io_out[9]
port 145 nsew signal output
rlabel metal3 s 104600 41328 105000 41384 6 irq[0]
port 146 nsew signal output
rlabel metal3 s 104600 42000 105000 42056 6 irq[1]
port 147 nsew signal output
rlabel metal3 s 104600 42672 105000 42728 6 irq[2]
port 148 nsew signal output
rlabel metal2 s 26208 69600 26264 70000 6 irqs[0]
port 149 nsew signal input
rlabel metal2 s 27552 69600 27608 70000 6 irqs[1]
port 150 nsew signal input
rlabel metal2 s 28896 69600 28952 70000 6 irqs[2]
port 151 nsew signal input
rlabel metal2 s 30240 69600 30296 70000 6 irqs[3]
port 152 nsew signal input
rlabel metal2 s 31584 69600 31640 70000 6 irqs[4]
port 153 nsew signal input
rlabel metal2 s 32928 69600 32984 70000 6 irqs[5]
port 154 nsew signal input
rlabel metal2 s 34272 69600 34328 70000 6 irqs[6]
port 155 nsew signal input
rlabel metal3 s 104600 3696 105000 3752 6 la_data_out[0]
port 156 nsew signal output
rlabel metal3 s 104600 10416 105000 10472 6 la_data_out[10]
port 157 nsew signal output
rlabel metal3 s 104600 11088 105000 11144 6 la_data_out[11]
port 158 nsew signal output
rlabel metal3 s 104600 11760 105000 11816 6 la_data_out[12]
port 159 nsew signal output
rlabel metal3 s 104600 12432 105000 12488 6 la_data_out[13]
port 160 nsew signal output
rlabel metal3 s 104600 13104 105000 13160 6 la_data_out[14]
port 161 nsew signal output
rlabel metal3 s 104600 13776 105000 13832 6 la_data_out[15]
port 162 nsew signal output
rlabel metal3 s 104600 14448 105000 14504 6 la_data_out[16]
port 163 nsew signal output
rlabel metal3 s 104600 15120 105000 15176 6 la_data_out[17]
port 164 nsew signal output
rlabel metal3 s 104600 15792 105000 15848 6 la_data_out[18]
port 165 nsew signal output
rlabel metal3 s 104600 16464 105000 16520 6 la_data_out[19]
port 166 nsew signal output
rlabel metal3 s 104600 4368 105000 4424 6 la_data_out[1]
port 167 nsew signal output
rlabel metal3 s 104600 17136 105000 17192 6 la_data_out[20]
port 168 nsew signal output
rlabel metal3 s 104600 17808 105000 17864 6 la_data_out[21]
port 169 nsew signal output
rlabel metal3 s 104600 18480 105000 18536 6 la_data_out[22]
port 170 nsew signal output
rlabel metal3 s 104600 19152 105000 19208 6 la_data_out[23]
port 171 nsew signal output
rlabel metal3 s 104600 19824 105000 19880 6 la_data_out[24]
port 172 nsew signal output
rlabel metal3 s 104600 20496 105000 20552 6 la_data_out[25]
port 173 nsew signal output
rlabel metal3 s 104600 21168 105000 21224 6 la_data_out[26]
port 174 nsew signal output
rlabel metal3 s 104600 21840 105000 21896 6 la_data_out[27]
port 175 nsew signal output
rlabel metal3 s 104600 22512 105000 22568 6 la_data_out[28]
port 176 nsew signal output
rlabel metal3 s 104600 23184 105000 23240 6 la_data_out[29]
port 177 nsew signal output
rlabel metal3 s 104600 5040 105000 5096 6 la_data_out[2]
port 178 nsew signal output
rlabel metal3 s 104600 23856 105000 23912 6 la_data_out[30]
port 179 nsew signal output
rlabel metal3 s 104600 24528 105000 24584 6 la_data_out[31]
port 180 nsew signal output
rlabel metal3 s 104600 25200 105000 25256 6 la_data_out[32]
port 181 nsew signal output
rlabel metal3 s 104600 25872 105000 25928 6 la_data_out[33]
port 182 nsew signal output
rlabel metal3 s 104600 26544 105000 26600 6 la_data_out[34]
port 183 nsew signal output
rlabel metal3 s 104600 27216 105000 27272 6 la_data_out[35]
port 184 nsew signal output
rlabel metal3 s 104600 27888 105000 27944 6 la_data_out[36]
port 185 nsew signal output
rlabel metal3 s 104600 28560 105000 28616 6 la_data_out[37]
port 186 nsew signal output
rlabel metal3 s 104600 29232 105000 29288 6 la_data_out[38]
port 187 nsew signal output
rlabel metal3 s 104600 29904 105000 29960 6 la_data_out[39]
port 188 nsew signal output
rlabel metal3 s 104600 5712 105000 5768 6 la_data_out[3]
port 189 nsew signal output
rlabel metal3 s 104600 30576 105000 30632 6 la_data_out[40]
port 190 nsew signal output
rlabel metal3 s 104600 31248 105000 31304 6 la_data_out[41]
port 191 nsew signal output
rlabel metal3 s 104600 31920 105000 31976 6 la_data_out[42]
port 192 nsew signal output
rlabel metal3 s 104600 32592 105000 32648 6 la_data_out[43]
port 193 nsew signal output
rlabel metal3 s 104600 33264 105000 33320 6 la_data_out[44]
port 194 nsew signal output
rlabel metal3 s 104600 33936 105000 33992 6 la_data_out[45]
port 195 nsew signal output
rlabel metal3 s 104600 34608 105000 34664 6 la_data_out[46]
port 196 nsew signal output
rlabel metal3 s 104600 35280 105000 35336 6 la_data_out[47]
port 197 nsew signal output
rlabel metal3 s 104600 35952 105000 36008 6 la_data_out[48]
port 198 nsew signal output
rlabel metal3 s 104600 36624 105000 36680 6 la_data_out[49]
port 199 nsew signal output
rlabel metal3 s 104600 6384 105000 6440 6 la_data_out[4]
port 200 nsew signal output
rlabel metal3 s 104600 37296 105000 37352 6 la_data_out[50]
port 201 nsew signal output
rlabel metal3 s 104600 37968 105000 38024 6 la_data_out[51]
port 202 nsew signal output
rlabel metal3 s 104600 38640 105000 38696 6 la_data_out[52]
port 203 nsew signal output
rlabel metal3 s 104600 39312 105000 39368 6 la_data_out[53]
port 204 nsew signal output
rlabel metal3 s 104600 39984 105000 40040 6 la_data_out[54]
port 205 nsew signal output
rlabel metal3 s 104600 40656 105000 40712 6 la_data_out[55]
port 206 nsew signal output
rlabel metal3 s 104600 7056 105000 7112 6 la_data_out[5]
port 207 nsew signal output
rlabel metal3 s 104600 7728 105000 7784 6 la_data_out[6]
port 208 nsew signal output
rlabel metal3 s 104600 8400 105000 8456 6 la_data_out[7]
port 209 nsew signal output
rlabel metal3 s 104600 9072 105000 9128 6 la_data_out[8]
port 210 nsew signal output
rlabel metal3 s 104600 9744 105000 9800 6 la_data_out[9]
port 211 nsew signal output
rlabel metal2 s 70560 69600 70616 70000 6 last_addr[0]
port 212 nsew signal output
rlabel metal2 s 84000 69600 84056 70000 6 last_addr[10]
port 213 nsew signal output
rlabel metal2 s 85344 69600 85400 70000 6 last_addr[11]
port 214 nsew signal output
rlabel metal2 s 86688 69600 86744 70000 6 last_addr[12]
port 215 nsew signal output
rlabel metal2 s 88032 69600 88088 70000 6 last_addr[13]
port 216 nsew signal output
rlabel metal2 s 89376 69600 89432 70000 6 last_addr[14]
port 217 nsew signal output
rlabel metal2 s 90720 69600 90776 70000 6 last_addr[15]
port 218 nsew signal output
rlabel metal2 s 71904 69600 71960 70000 6 last_addr[1]
port 219 nsew signal output
rlabel metal2 s 73248 69600 73304 70000 6 last_addr[2]
port 220 nsew signal output
rlabel metal2 s 74592 69600 74648 70000 6 last_addr[3]
port 221 nsew signal output
rlabel metal2 s 75936 69600 75992 70000 6 last_addr[4]
port 222 nsew signal output
rlabel metal2 s 77280 69600 77336 70000 6 last_addr[5]
port 223 nsew signal output
rlabel metal2 s 78624 69600 78680 70000 6 last_addr[6]
port 224 nsew signal output
rlabel metal2 s 79968 69600 80024 70000 6 last_addr[7]
port 225 nsew signal output
rlabel metal2 s 81312 69600 81368 70000 6 last_addr[8]
port 226 nsew signal output
rlabel metal2 s 82656 69600 82712 70000 6 last_addr[9]
port 227 nsew signal output
rlabel metal2 s 69216 69600 69272 70000 6 le_hi_act
port 228 nsew signal output
rlabel metal2 s 67872 69600 67928 70000 6 le_lo_act
port 229 nsew signal output
rlabel metal3 s 0 62496 400 62552 6 ram_bus_in[0]
port 230 nsew signal input
rlabel metal3 s 0 63168 400 63224 6 ram_bus_in[1]
port 231 nsew signal input
rlabel metal3 s 0 63840 400 63896 6 ram_bus_in[2]
port 232 nsew signal input
rlabel metal3 s 0 64512 400 64568 6 ram_bus_in[3]
port 233 nsew signal input
rlabel metal3 s 0 65184 400 65240 6 ram_bus_in[4]
port 234 nsew signal input
rlabel metal3 s 0 65856 400 65912 6 ram_bus_in[5]
port 235 nsew signal input
rlabel metal3 s 0 66528 400 66584 6 ram_bus_in[6]
port 236 nsew signal input
rlabel metal3 s 0 67200 400 67256 6 ram_bus_in[7]
port 237 nsew signal input
rlabel metal3 s 0 67872 400 67928 6 ram_enabled
port 238 nsew signal output
rlabel metal3 s 104600 56112 105000 56168 6 requested_addr[0]
port 239 nsew signal output
rlabel metal3 s 104600 62832 105000 62888 6 requested_addr[10]
port 240 nsew signal output
rlabel metal3 s 104600 63504 105000 63560 6 requested_addr[11]
port 241 nsew signal output
rlabel metal3 s 104600 64176 105000 64232 6 requested_addr[12]
port 242 nsew signal output
rlabel metal3 s 104600 64848 105000 64904 6 requested_addr[13]
port 243 nsew signal output
rlabel metal3 s 104600 65520 105000 65576 6 requested_addr[14]
port 244 nsew signal output
rlabel metal3 s 104600 66192 105000 66248 6 requested_addr[15]
port 245 nsew signal output
rlabel metal3 s 104600 56784 105000 56840 6 requested_addr[1]
port 246 nsew signal output
rlabel metal3 s 104600 57456 105000 57512 6 requested_addr[2]
port 247 nsew signal output
rlabel metal3 s 104600 58128 105000 58184 6 requested_addr[3]
port 248 nsew signal output
rlabel metal3 s 104600 58800 105000 58856 6 requested_addr[4]
port 249 nsew signal output
rlabel metal3 s 104600 59472 105000 59528 6 requested_addr[5]
port 250 nsew signal output
rlabel metal3 s 104600 60144 105000 60200 6 requested_addr[6]
port 251 nsew signal output
rlabel metal3 s 104600 60816 105000 60872 6 requested_addr[7]
port 252 nsew signal output
rlabel metal3 s 104600 61488 105000 61544 6 requested_addr[8]
port 253 nsew signal output
rlabel metal3 s 104600 62160 105000 62216 6 requested_addr[9]
port 254 nsew signal output
rlabel metal3 s 104600 49392 105000 49448 6 reset_out
port 255 nsew signal output
rlabel metal3 s 0 57120 400 57176 6 rom_bus_in[0]
port 256 nsew signal input
rlabel metal3 s 0 57792 400 57848 6 rom_bus_in[1]
port 257 nsew signal input
rlabel metal3 s 0 58464 400 58520 6 rom_bus_in[2]
port 258 nsew signal input
rlabel metal3 s 0 59136 400 59192 6 rom_bus_in[3]
port 259 nsew signal input
rlabel metal3 s 0 59808 400 59864 6 rom_bus_in[4]
port 260 nsew signal input
rlabel metal3 s 0 60480 400 60536 6 rom_bus_in[5]
port 261 nsew signal input
rlabel metal3 s 0 61152 400 61208 6 rom_bus_in[6]
port 262 nsew signal input
rlabel metal3 s 0 61824 400 61880 6 rom_bus_in[7]
port 263 nsew signal input
rlabel metal3 s 0 51744 400 51800 6 rom_bus_out[0]
port 264 nsew signal output
rlabel metal3 s 0 52416 400 52472 6 rom_bus_out[1]
port 265 nsew signal output
rlabel metal3 s 0 53088 400 53144 6 rom_bus_out[2]
port 266 nsew signal output
rlabel metal3 s 0 53760 400 53816 6 rom_bus_out[3]
port 267 nsew signal output
rlabel metal3 s 0 54432 400 54488 6 rom_bus_out[4]
port 268 nsew signal output
rlabel metal3 s 0 55104 400 55160 6 rom_bus_out[5]
port 269 nsew signal output
rlabel metal3 s 0 55776 400 55832 6 rom_bus_out[6]
port 270 nsew signal output
rlabel metal3 s 0 56448 400 56504 6 rom_bus_out[7]
port 271 nsew signal output
rlabel metal4 s 2224 1538 2384 68238 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 68238 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 68238 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 68238 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 68238 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 68238 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 68238 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 68238 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 68238 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 68238 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 68238 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 68238 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 68238 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 68238 6 vss
port 273 nsew ground bidirectional
rlabel metal2 s 1568 0 1624 400 6 wb_clk_i
port 274 nsew signal input
rlabel metal2 s 2576 0 2632 400 6 wb_rst_i
port 275 nsew signal input
rlabel metal2 s 3584 0 3640 400 6 wbs_ack_o
port 276 nsew signal output
rlabel metal2 s 7616 0 7672 400 6 wbs_adr_i[0]
port 277 nsew signal input
rlabel metal2 s 37856 0 37912 400 6 wbs_adr_i[10]
port 278 nsew signal input
rlabel metal2 s 40880 0 40936 400 6 wbs_adr_i[11]
port 279 nsew signal input
rlabel metal2 s 43904 0 43960 400 6 wbs_adr_i[12]
port 280 nsew signal input
rlabel metal2 s 46928 0 46984 400 6 wbs_adr_i[13]
port 281 nsew signal input
rlabel metal2 s 49952 0 50008 400 6 wbs_adr_i[14]
port 282 nsew signal input
rlabel metal2 s 52976 0 53032 400 6 wbs_adr_i[15]
port 283 nsew signal input
rlabel metal2 s 56000 0 56056 400 6 wbs_adr_i[16]
port 284 nsew signal input
rlabel metal2 s 59024 0 59080 400 6 wbs_adr_i[17]
port 285 nsew signal input
rlabel metal2 s 62048 0 62104 400 6 wbs_adr_i[18]
port 286 nsew signal input
rlabel metal2 s 65072 0 65128 400 6 wbs_adr_i[19]
port 287 nsew signal input
rlabel metal2 s 10640 0 10696 400 6 wbs_adr_i[1]
port 288 nsew signal input
rlabel metal2 s 68096 0 68152 400 6 wbs_adr_i[20]
port 289 nsew signal input
rlabel metal2 s 71120 0 71176 400 6 wbs_adr_i[21]
port 290 nsew signal input
rlabel metal2 s 74144 0 74200 400 6 wbs_adr_i[22]
port 291 nsew signal input
rlabel metal2 s 77168 0 77224 400 6 wbs_adr_i[23]
port 292 nsew signal input
rlabel metal2 s 80192 0 80248 400 6 wbs_adr_i[24]
port 293 nsew signal input
rlabel metal2 s 83216 0 83272 400 6 wbs_adr_i[25]
port 294 nsew signal input
rlabel metal2 s 86240 0 86296 400 6 wbs_adr_i[26]
port 295 nsew signal input
rlabel metal2 s 89264 0 89320 400 6 wbs_adr_i[27]
port 296 nsew signal input
rlabel metal2 s 92288 0 92344 400 6 wbs_adr_i[28]
port 297 nsew signal input
rlabel metal2 s 95312 0 95368 400 6 wbs_adr_i[29]
port 298 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 wbs_adr_i[2]
port 299 nsew signal input
rlabel metal2 s 98336 0 98392 400 6 wbs_adr_i[30]
port 300 nsew signal input
rlabel metal2 s 101360 0 101416 400 6 wbs_adr_i[31]
port 301 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 wbs_adr_i[3]
port 302 nsew signal input
rlabel metal2 s 19712 0 19768 400 6 wbs_adr_i[4]
port 303 nsew signal input
rlabel metal2 s 22736 0 22792 400 6 wbs_adr_i[5]
port 304 nsew signal input
rlabel metal2 s 25760 0 25816 400 6 wbs_adr_i[6]
port 305 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 wbs_adr_i[7]
port 306 nsew signal input
rlabel metal2 s 31808 0 31864 400 6 wbs_adr_i[8]
port 307 nsew signal input
rlabel metal2 s 34832 0 34888 400 6 wbs_adr_i[9]
port 308 nsew signal input
rlabel metal2 s 4592 0 4648 400 6 wbs_cyc_i
port 309 nsew signal input
rlabel metal2 s 8624 0 8680 400 6 wbs_dat_i[0]
port 310 nsew signal input
rlabel metal2 s 38864 0 38920 400 6 wbs_dat_i[10]
port 311 nsew signal input
rlabel metal2 s 41888 0 41944 400 6 wbs_dat_i[11]
port 312 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 wbs_dat_i[12]
port 313 nsew signal input
rlabel metal2 s 47936 0 47992 400 6 wbs_dat_i[13]
port 314 nsew signal input
rlabel metal2 s 50960 0 51016 400 6 wbs_dat_i[14]
port 315 nsew signal input
rlabel metal2 s 53984 0 54040 400 6 wbs_dat_i[15]
port 316 nsew signal input
rlabel metal2 s 57008 0 57064 400 6 wbs_dat_i[16]
port 317 nsew signal input
rlabel metal2 s 60032 0 60088 400 6 wbs_dat_i[17]
port 318 nsew signal input
rlabel metal2 s 63056 0 63112 400 6 wbs_dat_i[18]
port 319 nsew signal input
rlabel metal2 s 66080 0 66136 400 6 wbs_dat_i[19]
port 320 nsew signal input
rlabel metal2 s 11648 0 11704 400 6 wbs_dat_i[1]
port 321 nsew signal input
rlabel metal2 s 69104 0 69160 400 6 wbs_dat_i[20]
port 322 nsew signal input
rlabel metal2 s 72128 0 72184 400 6 wbs_dat_i[21]
port 323 nsew signal input
rlabel metal2 s 75152 0 75208 400 6 wbs_dat_i[22]
port 324 nsew signal input
rlabel metal2 s 78176 0 78232 400 6 wbs_dat_i[23]
port 325 nsew signal input
rlabel metal2 s 81200 0 81256 400 6 wbs_dat_i[24]
port 326 nsew signal input
rlabel metal2 s 84224 0 84280 400 6 wbs_dat_i[25]
port 327 nsew signal input
rlabel metal2 s 87248 0 87304 400 6 wbs_dat_i[26]
port 328 nsew signal input
rlabel metal2 s 90272 0 90328 400 6 wbs_dat_i[27]
port 329 nsew signal input
rlabel metal2 s 93296 0 93352 400 6 wbs_dat_i[28]
port 330 nsew signal input
rlabel metal2 s 96320 0 96376 400 6 wbs_dat_i[29]
port 331 nsew signal input
rlabel metal2 s 14672 0 14728 400 6 wbs_dat_i[2]
port 332 nsew signal input
rlabel metal2 s 99344 0 99400 400 6 wbs_dat_i[30]
port 333 nsew signal input
rlabel metal2 s 102368 0 102424 400 6 wbs_dat_i[31]
port 334 nsew signal input
rlabel metal2 s 17696 0 17752 400 6 wbs_dat_i[3]
port 335 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 wbs_dat_i[4]
port 336 nsew signal input
rlabel metal2 s 23744 0 23800 400 6 wbs_dat_i[5]
port 337 nsew signal input
rlabel metal2 s 26768 0 26824 400 6 wbs_dat_i[6]
port 338 nsew signal input
rlabel metal2 s 29792 0 29848 400 6 wbs_dat_i[7]
port 339 nsew signal input
rlabel metal2 s 32816 0 32872 400 6 wbs_dat_i[8]
port 340 nsew signal input
rlabel metal2 s 35840 0 35896 400 6 wbs_dat_i[9]
port 341 nsew signal input
rlabel metal2 s 9632 0 9688 400 6 wbs_dat_o[0]
port 342 nsew signal output
rlabel metal2 s 39872 0 39928 400 6 wbs_dat_o[10]
port 343 nsew signal output
rlabel metal2 s 42896 0 42952 400 6 wbs_dat_o[11]
port 344 nsew signal output
rlabel metal2 s 45920 0 45976 400 6 wbs_dat_o[12]
port 345 nsew signal output
rlabel metal2 s 48944 0 49000 400 6 wbs_dat_o[13]
port 346 nsew signal output
rlabel metal2 s 51968 0 52024 400 6 wbs_dat_o[14]
port 347 nsew signal output
rlabel metal2 s 54992 0 55048 400 6 wbs_dat_o[15]
port 348 nsew signal output
rlabel metal2 s 58016 0 58072 400 6 wbs_dat_o[16]
port 349 nsew signal output
rlabel metal2 s 61040 0 61096 400 6 wbs_dat_o[17]
port 350 nsew signal output
rlabel metal2 s 64064 0 64120 400 6 wbs_dat_o[18]
port 351 nsew signal output
rlabel metal2 s 67088 0 67144 400 6 wbs_dat_o[19]
port 352 nsew signal output
rlabel metal2 s 12656 0 12712 400 6 wbs_dat_o[1]
port 353 nsew signal output
rlabel metal2 s 70112 0 70168 400 6 wbs_dat_o[20]
port 354 nsew signal output
rlabel metal2 s 73136 0 73192 400 6 wbs_dat_o[21]
port 355 nsew signal output
rlabel metal2 s 76160 0 76216 400 6 wbs_dat_o[22]
port 356 nsew signal output
rlabel metal2 s 79184 0 79240 400 6 wbs_dat_o[23]
port 357 nsew signal output
rlabel metal2 s 82208 0 82264 400 6 wbs_dat_o[24]
port 358 nsew signal output
rlabel metal2 s 85232 0 85288 400 6 wbs_dat_o[25]
port 359 nsew signal output
rlabel metal2 s 88256 0 88312 400 6 wbs_dat_o[26]
port 360 nsew signal output
rlabel metal2 s 91280 0 91336 400 6 wbs_dat_o[27]
port 361 nsew signal output
rlabel metal2 s 94304 0 94360 400 6 wbs_dat_o[28]
port 362 nsew signal output
rlabel metal2 s 97328 0 97384 400 6 wbs_dat_o[29]
port 363 nsew signal output
rlabel metal2 s 15680 0 15736 400 6 wbs_dat_o[2]
port 364 nsew signal output
rlabel metal2 s 100352 0 100408 400 6 wbs_dat_o[30]
port 365 nsew signal output
rlabel metal2 s 103376 0 103432 400 6 wbs_dat_o[31]
port 366 nsew signal output
rlabel metal2 s 18704 0 18760 400 6 wbs_dat_o[3]
port 367 nsew signal output
rlabel metal2 s 21728 0 21784 400 6 wbs_dat_o[4]
port 368 nsew signal output
rlabel metal2 s 24752 0 24808 400 6 wbs_dat_o[5]
port 369 nsew signal output
rlabel metal2 s 27776 0 27832 400 6 wbs_dat_o[6]
port 370 nsew signal output
rlabel metal2 s 30800 0 30856 400 6 wbs_dat_o[7]
port 371 nsew signal output
rlabel metal2 s 33824 0 33880 400 6 wbs_dat_o[8]
port 372 nsew signal output
rlabel metal2 s 36848 0 36904 400 6 wbs_dat_o[9]
port 373 nsew signal output
rlabel metal2 s 5600 0 5656 400 6 wbs_stb_i
port 374 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 wbs_we_i
port 375 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 105000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 14822628
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/AS2650/openlane/wrapped_as2650/runs/23_11_27_22_59/results/signoff/wrapped_as2650.magic.gds
string GDS_START 581818
<< end >>

